`timescale 1 ns/100 ps
// Version: v11.8 SP3 11.8.3.6


module sig_gen_9(
       inc_const_c,
       n_rst_c,
       clk_c,
       inc_constd
    );
input  inc_const_c;
input  n_rst_c;
input  clk_c;
output inc_constd;

    wire sig_prev_i, sig_prev_net_1, sig_old_i_0, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(clk_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev (.D(inc_const_c), .CLK(clk_c), .CLR(n_rst_c), .Q(
        sig_prev_net_1));
    INV sig_old_RNO (.A(sig_prev_net_1), .Y(sig_prev_i));
    NOR2B sig_old_RNIK1HQ (.A(sig_old_i_0), .B(sig_prev_net_1), .Y(
        inc_constd));
    GND GND_i (.Y(GND));
    
endmodule


module pwm_ctl_400s_32s_13s_0_1_2_3(
       sum_8,
       sum_39,
       sum_9,
       sum_10,
       sum_11,
       sum_12,
       sum_13,
       sum_14,
       sum_16,
       sum_18,
       sum_19,
       sum_20,
       sum_21,
       sum_23,
       sum_22,
       sum_17,
       sum_15,
       sum_1_d0,
       sum_0_d0,
       sum_2_d0,
       sum_7,
       sum_6,
       sum_4,
       sum_3,
       sum_5,
       off_div,
       sum_2_0,
       sum_1_0,
       sum_0_0,
       state,
       n_rst_c,
       clk_c,
       pwm_enable
    );
input  sum_8;
input  sum_39;
input  sum_9;
input  sum_10;
input  sum_11;
input  sum_12;
input  sum_13;
input  sum_14;
input  sum_16;
input  sum_18;
input  sum_19;
input  sum_20;
input  sum_21;
input  sum_23;
input  sum_22;
input  sum_17;
input  sum_15;
input  sum_1_d0;
input  sum_0_d0;
input  sum_2_d0;
input  sum_7;
input  sum_6;
input  sum_4;
input  sum_3;
input  sum_5;
output [31:0] off_div;
input  sum_2_0;
input  sum_1_0;
input  sum_0_0;
output [1:0] state;
input  n_rst_c;
input  clk_c;
input  pwm_enable;

    wire \state_d_0[2] , un1_state_2_0, un5lt31, 
        next_off_div_2_sqmuxa_11, N_16, \DWACT_FINC_E[4] , N_13, 
        \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , ADD_32x32_fast_I321_Y_0, 
        ADD_32x32_fast_I258_Y_3, N610, N625, ADD_32x32_fast_I258_Y_2, 
        N482, ADD_32x32_fast_I258_Y_0, N551, ADD_32x32_fast_I320_Y_0, 
        ADD_32x32_fast_I313_Y_0, ADD_32x32_fast_I259_Y_3, N612, N627, 
        ADD_32x32_fast_I259_Y_2, N484, ADD_32x32_fast_I259_Y_0, N553, 
        ADD_32x32_fast_I258_un1_Y_0, N626, ADD_32x32_fast_I318_Y_0, 
        ADD_32x32_fast_I319_Y_0, ADD_32x32_fast_I317_Y_0, 
        ADD_32x32_fast_I314_Y_0, ADD_32x32_fast_I316_Y_0, 
        ADD_32x32_fast_I315_Y_0, ADD_32x32_fast_I266_Y_0, N641, 
        ADD_32x32_fast_I260_Y_2, N614, N629, ADD_32x32_fast_I260_Y_1, 
        N486, N555, ADD_32x32_fast_I261_Y_2, N616, N631, 
        ADD_32x32_fast_I261_Y_1, N488, N557, ADD_32x32_fast_I312_Y_0, 
        ADD_32x32_fast_I304_Y_0, \un1_sum_adj[14] , 
        ADD_32x32_fast_I259_un1_Y_0, N628, ADD_32x32_fast_I262_Y_1, 
        N618, N633, ADD_32x32_fast_I262_Y_0, N559, 
        ADD_32x32_fast_I310_Y_0, ADD_32x32_fast_I311_Y_0, 
        ADD_32x32_fast_I309_Y_0, ADD_32x32_fast_I266_un1_Y_0, N642, 
        ADD_32x32_fast_I265_Y_0, N565, ADD_32x32_fast_I264_Y_1, N622, 
        N637, ADD_32x32_fast_I264_Y_0, N563, ADD_32x32_fast_I263_Y_1, 
        N620, N635, ADD_32x32_fast_I263_Y_0, N561, 
        ADD_32x32_fast_I308_Y_0, ADD_32x32_fast_I307_Y_0, 
        ADD_32x32_fast_I306_Y_0, ADD_32x32_fast_I303_Y_0, 
        \sum_adj[21]_net_1 , ADD_32x32_fast_I302_Y_0, 
        \un1_sum_adj[12] , ADD_32x32_fast_I261_un1_Y_0, N632, 
        ADD_32x32_fast_I260_un1_Y_0, N630, ADD_32x32_fast_I301_Y_0, 
        \sum_adj[19]_net_1 , ADD_32x32_fast_I262_un1_Y_0, N634, 
        ADD_32x32_fast_I269_Y_0, N647, ADD_32x32_fast_I270_Y_0, N649, 
        ADD_32x32_fast_I299_Y_0, \sum_adj[17]_net_1 , 
        ADD_32x32_fast_I300_Y_0, \un1_sum_adj[10] , 
        ADD_32x32_fast_I298_Y_0, \un1_sum_adj[8] , 
        ADD_32x32_fast_I263_un1_Y_0, N636, ADD_32x32_fast_I264_un1_Y_0, 
        N638, ADD_32x32_fast_I265_un1_Y_0, N624, N640, 
        ADD_32x32_fast_I296_Y_0, \sum_adj[14]_net_1 , 
        ADD_32x32_fast_I271_Y_0, ADD_32x32_fast_I271_un1_Y_0, 
        ADD_32x32_fast_I273_Y_0, ADD_32x32_fast_I273_un1_Y_0, N639, 
        ADD_32x32_fast_I272_Y_0, ADD_32x32_fast_I272_un1_Y_0, 
        ADD_32x32_fast_I295_Y_0, \un1_sum_adj[5] , 
        ADD_32x32_fast_I294_Y_0, \sum_adj[12]_net_1 , 
        ADD_32x32_fast_I293_Y_0, \un1_sum_adj[3] , N538, N654, N590, 
        N598, \un1_sum_adj[0] , N586, N594, N601, 
        ADD_32x32_fast_I292_Y_0, \sum_adj[10]_net_1 , 
        next_off_div_2_sqmuxa_9, next_off_div_2_sqmuxa_8, 
        next_off_div37, next_off_div_2_sqmuxa_1, 
        next_off_div_2_sqmuxa_0, next_off_div_2_sqmuxa_7, 
        un1_off_divlto31_10, next_off_div_2_sqmuxa_5, 
        next_off_div_2_sqmuxa_3, ADD_32x32_fast_I291_Y_0, 
        \un1_sum_adj[1] , un5lto20_2, un5lto20_1, 
        ADD_32x32_fast_I155_Y_0, ADD_32x32_fast_I157_Y_0, un5lto14_2, 
        un5lto14_1, un1_off_divlto31_22, un1_off_divlto31_15, 
        un1_off_divlto31_14, un1_off_divlto31_20, un1_off_divlto31_21, 
        un1_off_divlto31_13, un1_off_divlto31_12, un1_off_divlto31_17, 
        un1_off_divlto31_9, un1_off_divlt31, un1_off_divlto31_0, 
        un5lto9, un1_off_divlto31_8, un1_off_divlto31_6, 
        un1_off_divlto31_4, un1_off_divlto31_2, un5lto7_1, I269_un1_Y, 
        N648, N663, I270_un1_Y, N650, N599, \un1_off_div_1[7] , 
        \un1_sum_adj[7] , N657, \un1_off_div_1[20] , 
        \un1_off_div_1[19] , \un1_off_div_1[18] , I236_un1_Y, 
        \un1_off_div_1[10] , N796, N765, N779, N655, 
        \un1_off_div_1[15] , \un1_sum_adj[15] , N781, N485, N489, N558, 
        N755, N790, I262_un1_Y, N793, I265_un1_Y, N802, N763, 
        I224_un1_Y, \un1_off_div_1[27] , N759, N751, N784, N554, N753, 
        N787, N483, N487, N556, N552, N749, N761, N799, 
        \un1_off_div_1[17] , I238_un1_Y, un5lt16, I268_un1_Y, N646, 
        N661, N769, I230_un1_Y, un5lt9, un5lto4, un5lt4, 
        \un1_off_div_1[5] , \un1_off_div_1[0] , \un1_off_div_1[3] , 
        N767, I228_un1_Y, I267_un1_Y, N644, N659, \nsum_adj_11[8] , 
        I_23_5, \nsum_adj_11[9] , I_26_1, \nsum_adj_11[10] , I_28_1, 
        \nsum_adj_11[11] , I_32_1, \nsum_adj_11[12] , I_35_1, 
        \nsum_adj_11[13] , I_37_1, \nsum_adj_11[14] , I_40_1, 
        \nsum_adj_11[16] , I_46_1, \nsum_adj_11[18] , I_53_1, 
        \nsum_adj_11[19] , I_56_1, \nsum_adj_11[20] , I_59_1, 
        \nsum_adj_11[21] , I_62_1, \nsum_adj_11[23] , I_70_1, 
        \state_ns[0] , state_176_d, \nsum_adj_11[22] , I_65_1, N_311_i, 
        \nsum_adj_11[17] , I_49_1, \nsum_adj_11[15] , I_43_1, 
        \next_off_div[1] , \next_off_div[2] , \next_off_div[8] , 
        \next_off_div[9] , \next_off_div[11] , \next_off_div[12] , 
        \next_off_div[22] , \state_d[2] , N383, N386, N387, N390, N392, 
        N395, N396, N404, N408, N521, N411, N522, N407, N523, N528, 
        N529, N530, N531, N532, N389, N533, N534, N535, N536, N537, 
        \sum_adj[8]_net_1 , N525, N589, N524, N593, N595, N596, N597, 
        I150_un1_Y, N564, N572, N579, N571, N580, N645, N587, N588, 
        N653, I204_un1_Y, N518, N515, N514, N416, N420, N419, N417, 
        N576, N511, N507, N510, N506, N519, N413, N513, N423, N516, 
        N517, N410, N520, N575, N578, N581, N582, N585, N643, 
        I246_un1_Y, \sum_adj[20]_net_1 , \sum_adj[18]_net_1 , 
        \sum_adj[16]_net_1 , \sum_adj[15]_net_1 , \sum_adj[11]_net_1 , 
        \sum_adj[9]_net_1 , \next_off_div[3] , next_off_div_0_sqmuxa, 
        \next_off_div[0] , \next_off_div[5] , N591, N584, N583, N568, 
        N567, N560, N503, N502, N592, N527, N402, N401, N426, N432, 
        N428, N429, \sum_adj[13]_net_1 , N398, \next_off_div[21] , 
        N577, \next_off_div[14] , next_off_div_1_sqmuxa, un1_state_2, 
        un5lt14, \next_off_div[17] , \next_off_div[31] , 
        \next_off_div[25] , N490, N491, N494, \next_off_div[29] , 
        \next_off_div[30] , N562, N492, N493, N496, N566, N573, 
        \next_off_div[26] , I249_un1_Y, N574, I184_un1_Y, N509, 
        \next_off_div[28] , \next_off_div[27] , \next_off_div[24] , 
        N495, N497, N425, N508, N422, \sum_adj[23]_net_1 , 
        \sum_adj[22]_net_1 , \next_off_div[15] , \next_off_div[6] , 
        N526, N498, N499, N512, \next_off_div[13] , \next_off_div[16] , 
        N569, N570, N500, N501, N504, N505, \next_off_div[23] , 
        \next_off_div[7] , \next_off_div[10] , \next_off_div[18] , 
        \next_off_div[19] , \next_off_div[20] , I247_un1_Y, N651, 
        I196_un1_Y, \next_off_div[4] , N_2, \DWACT_FINC_E[29] , 
        \DWACT_FINC_E[13] , \DWACT_FINC_E[33] , \DWACT_FINC_E[34] , 
        \DWACT_FINC_E[2] , \DWACT_FINC_E[5] , \DWACT_FINC_E[15] , N_3, 
        \DWACT_FINC_E[28] , \DWACT_FINC_E[16] , N_4, N_5, 
        \DWACT_FINC_E[14] , N_6, \DWACT_FINC_E[9] , \DWACT_FINC_E[12] , 
        N_7, \DWACT_FINC_E[10] , \DWACT_FINC_E[0] , N_8, 
        \DWACT_FINC_E[11] , N_9, N_10, N_11, \DWACT_FINC_E[8] , N_12, 
        N_14, N_15, \DWACT_FINC_E[3] , N_17, GND, VCC;
    
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I59_Y (.A(sum_1_0), .B(
        off_div[17]), .C(N432), .Y(N505));
    AO1 \off_div_RNIOMI84[31]  (.A(un1_off_divlto31_22), .B(
        un1_off_divlto31_21), .C(off_div[31]), .Y(next_off_div37));
    NOR2B \off_div_RNI2MK4[19]  (.A(off_div[20]), .B(off_div[19]), .Y(
        un5lto20_1));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_2 (.A(N482), .B(
        ADD_32x32_fast_I258_Y_0), .C(N551), .Y(ADD_32x32_fast_I258_Y_2)
        );
    DFN1C0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(state[0]));
    DFN1E0C0 \off_div[29]  (.D(\next_off_div[29] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[29]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y_0 (.A(N555), .B(N563), 
        .Y(ADD_32x32_fast_I264_Y_0));
    DFN1E0C0 \off_div[26]  (.D(\next_off_div[26] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[26]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I247_Y (.A(I247_un1_Y), .B(
        N651), .Y(N796));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I108_Y (.A(N496), .B(N492), 
        .Y(N557));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I47_Y (.A(off_div[23]), .B(
        off_div[22]), .C(sum_0_0), .Y(N493));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I165_Y (.A(N562), .B(N554), 
        .Y(N620));
    XNOR2 un13_nsum_adj_I_49 (.A(sum_17), .B(N_8), .Y(I_49_1));
    NOR3 un13_nsum_adj_I_10 (.A(sum_1_d0), .B(sum_0_d0), .C(sum_2_d0), 
        .Y(\DWACT_FINC_E[0] ));
    DFN1E0C0 \off_div[31]  (.D(\next_off_div[31] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[31]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I149_Y (.A(N537), .B(N533), 
        .Y(N598));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I135_Y (.A(N519), .B(N523), 
        .Y(N584));
    AND3 un13_nsum_adj_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[6] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I147_Y (.A(N535), .B(N531), 
        .Y(N596));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I121_Y (.A(N505), .B(N509), 
        .Y(N570));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I272_Y_0 (.A(
        ADD_32x32_fast_I272_un1_Y_0), .B(N638), .C(N637), .Y(
        ADD_32x32_fast_I272_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I173_Y (.A(N562), .B(N570), 
        .Y(N628));
    MX2 \sum_adj_RNO[9]  (.A(sum_9), .B(I_26_1), .S(sum_2_0), .Y(
        \nsum_adj_11[9] ));
    XA1 \off_div_RNO[22]  (.A(N767), .B(ADD_32x32_fast_I312_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[22] ));
    DFN1E1C0 \sum_adj[23]  (.D(\nsum_adj_11[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[23]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I203_Y (.A(N594), .B(N601), 
        .C(N593), .Y(N659));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I155_Y (.A(N483), .B(
        ADD_32x32_fast_I155_Y_0), .C(N552), .Y(N610));
    NOR2 un13_nsum_adj_I_57 (.A(sum_18), .B(sum_19), .Y(
        \DWACT_FINC_E[14] ));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I86_Y (.A(N389), .B(
        off_div[3]), .C(\un1_sum_adj[3] ), .Y(N532));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I200_Y (.A(N597), .B(N590), 
        .C(N589), .Y(N655));
    MX2 \sum_adj_RNO[15]  (.A(sum_15), .B(I_43_1), .S(sum_1_0), .Y(
        \nsum_adj_11[15] ));
    XNOR2 un13_nsum_adj_I_53 (.A(sum_18), .B(N_7), .Y(I_53_1));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I315_Y_0 (.A(off_div[25]), 
        .B(sum_39), .Y(ADD_32x32_fast_I315_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I84_Y (.A(N392), .B(N396), .C(
        N395), .Y(N530));
    NOR3B un13_nsum_adj_I_45 (.A(\DWACT_FINC_E[10] ), .B(
        \DWACT_FINC_E[6] ), .C(sum_15), .Y(N_9));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I130_Y (.A(N518), .B(N515), 
        .C(N514), .Y(N579));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I266_Y (.A(
        ADD_32x32_fast_I266_un1_Y_0), .B(N657), .C(
        ADD_32x32_fast_I266_Y_0), .Y(N765));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I118_Y (.A(N506), .B(N503), 
        .C(N502), .Y(N567));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I273_un1_Y_0 (.A(N590), .B(
        N598), .C(\un1_sum_adj[0] ), .Y(ADD_32x32_fast_I273_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I69_Y (.A(N417), .B(N420), 
        .Y(N515));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I262_Y_0 (.A(N551), .B(N559), 
        .Y(ADD_32x32_fast_I262_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I202_Y (.A(N592), .B(N599), 
        .C(N591), .Y(N657));
    OR2 \off_div_RNI7PCO[8]  (.A(off_div[9]), .B(off_div[8]), .Y(
        un5lto9));
    MX2 \sum_adj_RNO[16]  (.A(sum_16), .B(I_46_1), .S(sum_1_0), .Y(
        \nsum_adj_11[16] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I309_Y_0 (.A(off_div[19]), 
        .B(sum_39), .Y(ADD_32x32_fast_I309_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I184_un1_Y (.A(N581), .B(
        N574), .Y(I184_un1_Y));
    MX2 \off_div_RNO[3]  (.A(next_off_div_0_sqmuxa), .B(
        \un1_off_div_1[3] ), .S(\state_d_0[2] ), .Y(\next_off_div[3] ));
    AND3 un13_nsum_adj_I_69 (.A(\DWACT_FINC_E[29] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[33] ), .Y(N_2));
    AO1C \state_RNI3P9DA_0[1]  (.A(un5lt31), .B(
        next_off_div_2_sqmuxa_11), .C(state[1]), .Y(un1_state_2_0));
    OA1 \off_div_RNI7A8S3[10]  (.A(un5lto9), .B(un5lt9), .C(
        off_div[10]), .Y(un5lt14));
    OA1 \off_div_RNIKRH13[1]  (.A(un5lto4), .B(un5lt4), .C(un5lto7_1), 
        .Y(un5lt9));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I76_Y (.A(N404), .B(N408), .C(
        N407), .Y(N522));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I4_G0N (.A(sum_0_0), .B(
        \sum_adj[12]_net_1 ), .C(off_div[4]), .Y(N395));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I1_P0N (.A(\un1_sum_adj[1] ), 
        .B(off_div[1]), .Y(N387));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I13_G0N (.A(sum_2_0), .B(
        \sum_adj[21]_net_1 ), .C(off_div[13]), .Y(N422));
    DFN1E0C0 \off_div[15]  (.D(\next_off_div[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[15]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I150_Y (.A(I150_un1_Y), .B(
        N534), .Y(N599));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I144_Y (.A(N532), .B(N529), 
        .C(N528), .Y(N593));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I74_Y (.A(N407), .B(N411), .C(
        N410), .Y(N520));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I50_Y (.A(off_div[20]), .B(
        off_div[21]), .C(sum_0_0), .Y(N496));
    DFN1E0C0 \off_div[13]  (.D(\next_off_div[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[13]));
    MX2 \sum_adj_RNO[20]  (.A(sum_20), .B(I_59_1), .S(sum_1_0), .Y(
        \nsum_adj_11[20] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I293_Y_0 (.A(off_div[3]), .B(
        \un1_sum_adj[3] ), .Y(ADD_32x32_fast_I293_Y_0));
    AND2 un13_nsum_adj_I_44 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[9] ), .Y(\DWACT_FINC_E[10] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I272_un1_Y_0 (.A(N538), .B(
        N654), .Y(ADD_32x32_fast_I272_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I265_un1_Y (.A(
        ADD_32x32_fast_I265_un1_Y_0), .B(N802), .Y(I265_un1_Y));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I319_Y_0 (.A(off_div[29]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I319_Y_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I265_Y_0 (.A(N557), .B(N565), 
        .Y(ADD_32x32_fast_I265_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I179_Y (.A(N576), .B(N568), 
        .Y(N634));
    AND3 un13_nsum_adj_I_39 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[8] ), .Y(N_11));
    XA1 \off_div_RNO[24]  (.A(N763), .B(ADD_32x32_fast_I314_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[24] ));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I309_Y (.A(I270_un1_Y), .B(
        ADD_32x32_fast_I270_Y_0), .C(ADD_32x32_fast_I309_Y_0), .Y(
        \un1_off_div_1[19] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I177_Y (.A(N566), .B(N574), 
        .Y(N632));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I51_Y (.A(off_div[21]), .B(
        off_div[20]), .C(sum_0_0), .Y(N497));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I308_Y_0 (.A(off_div[18]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I308_Y_0));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I2_P0N (.A(sum_2_0), .B(
        \sum_adj[10]_net_1 ), .C(off_div[2]), .Y(N390));
    DFN1E0P0 \off_div[7]  (.D(\next_off_div[7] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2), .Q(off_div[7]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I196_Y (.A(I196_un1_Y), .B(
        N585), .Y(N651));
    NOR3 un13_nsum_adj_I_29 (.A(sum_7), .B(sum_6), .C(sum_8), .Y(
        \DWACT_FINC_E[5] ));
    XNOR2 un13_nsum_adj_I_65 (.A(sum_22), .B(N_3), .Y(I_65_1));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I268_Y (.A(I230_un1_Y), .B(
        N629), .C(I268_un1_Y), .Y(N769));
    DFN1E0C0 \off_div[9]  (.D(\next_off_div[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[9]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I37_Y (.A(off_div[28]), .B(
        off_div[27]), .C(sum_0_0), .Y(N483));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I186_Y (.A(N583), .B(N576), 
        .C(N575), .Y(N641));
    DFN1E0C0 \off_div[11]  (.D(\next_off_div[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[11]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I145_Y (.A(N533), .B(N529), 
        .Y(N594));
    DFN1E1C0 \sum_adj[18]  (.D(\nsum_adj_11[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[18]_net_1 ));
    MX2 un1_off_div_1_0_0_ADD_32x32_fast_I92_Y (.A(sum_2_0), .B(
        off_div[0]), .S(\sum_adj[8]_net_1 ), .Y(N538));
    XA1 \off_div_RNO[13]  (.A(N787), .B(ADD_32x32_fast_I303_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[13] ));
    NOR3C \off_div_RNI3UI41[6]  (.A(off_div[5]), .B(off_div[7]), .C(
        off_div[6]), .Y(un5lto7_1));
    MX2 \sum_adj_RNO[21]  (.A(sum_21), .B(I_62_1), .S(sum_1_0), .Y(
        \nsum_adj_11[21] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I318_Y_0 (.A(off_div[28]), 
        .B(sum_39), .Y(ADD_32x32_fast_I318_Y_0));
    XNOR2 un13_nsum_adj_I_35 (.A(sum_12), .B(N_13), .Y(I_35_1));
    XOR2 \sum_adj_RNILP5T[8]  (.A(\sum_adj[8]_net_1 ), .B(sum_39), .Y(
        \un1_sum_adj[0] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I191_Y (.A(N580), .B(N588), 
        .Y(N646));
    MX2 \sum_adj_RNO[22]  (.A(sum_22), .B(I_65_1), .S(sum_2_0), .Y(
        \nsum_adj_11[22] ));
    MX2 \off_div_RNO[15]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[15] ), .S(\state_d[2] ), .Y(\next_off_div[15] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y (.A(
        ADD_32x32_fast_I258_un1_Y_0), .B(N781), .C(
        ADD_32x32_fast_I258_Y_3), .Y(N749));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I14_P0N (.A(\un1_sum_adj[14] )
        , .B(off_div[14]), .Y(N426));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I122_Y (.A(N510), .B(N507), 
        .C(N506), .Y(N571));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I89_Y (.A(N387), .B(N390), 
        .Y(N535));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I262_Y_1 (.A(N618), .B(N633), 
        .C(ADD_32x32_fast_I262_Y_0), .Y(ADD_32x32_fast_I262_Y_1));
    AND3 un13_nsum_adj_I_64 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[16] ), .Y(N_3));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I265_Y (.A(I224_un1_Y), .B(
        ADD_32x32_fast_I265_Y_0), .C(I265_un1_Y), .Y(N763));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I181_Y (.A(N570), .B(N578), 
        .Y(N636));
    NOR2A un13_nsum_adj_I_25 (.A(\DWACT_FINC_E[4] ), .B(sum_8), .Y(
        N_16));
    DFN1E1C0 \sum_adj[9]  (.D(\nsum_adj_11[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[9]_net_1 ));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I60_Y (.A(N428), .B(sum_1_0), 
        .C(off_div[16]), .Y(N506));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I4_P0N (.A(sum_0_0), .B(
        \sum_adj[12]_net_1 ), .C(off_div[4]), .Y(N396));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I307_Y (.A(I238_un1_Y), .B(
        ADD_32x32_fast_I272_Y_0), .C(ADD_32x32_fast_I307_Y_0), .Y(
        \un1_off_div_1[17] ));
    AND3 un13_nsum_adj_I_51 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[28] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I174_Y (.A(N571), .B(N564), 
        .C(N563), .Y(N629));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I140_Y (.A(N528), .B(N525), 
        .C(N524), .Y(N589));
    DFN1E1C0 \sum_adj[11]  (.D(\nsum_adj_11[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[11]_net_1 ));
    NOR2A \off_div_RNIEO4E[31]  (.A(state[0]), .B(off_div[31]), .Y(
        next_off_div_2_sqmuxa_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y_1 (.A(N620), .B(N635), 
        .C(ADD_32x32_fast_I263_Y_0), .Y(ADD_32x32_fast_I263_Y_1));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I246_Y (.A(I246_un1_Y), .B(
        N649), .Y(N793));
    NOR2B \off_div_RNO[27]  (.A(\un1_off_div_1[27] ), .B(\state_d[2] ), 
        .Y(\next_off_div[27] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I291_Y_0 (.A(off_div[1]), .B(
        \un1_sum_adj[1] ), .Y(ADD_32x32_fast_I291_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I249_un1_Y (.A(N590), .B(
        N598), .C(\un1_sum_adj[0] ), .Y(I249_un1_Y));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I13_P0N (.A(sum_2_0), .B(
        \sum_adj[21]_net_1 ), .C(off_div[13]), .Y(N423));
    AND3 un13_nsum_adj_I_48 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[11] ), .Y(N_8));
    DFN1E0C0 \off_div[25]  (.D(\next_off_div[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[25]));
    XA1 \off_div_RNO[1]  (.A(N538), .B(ADD_32x32_fast_I291_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[1] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I61_Y (.A(N432), .B(N429), 
        .Y(N507));
    NOR2B un13_nsum_adj_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_13));
    DFN1E1C0 \sum_adj[22]  (.D(\nsum_adj_11[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[22]_net_1 ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I79_Y (.A(off_div[7]), .B(
        \un1_sum_adj[7] ), .C(N402), .Y(N525));
    OA1 \off_div_RNII4P74[15]  (.A(un5lt14), .B(un5lto14_2), .C(
        off_div[15]), .Y(un5lt16));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I150_un1_Y (.A(N535), .B(
        N538), .Y(I150_un1_Y));
    DFN1E0C0 \off_div[23]  (.D(\next_off_div[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[23]));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I304_Y_0 (.A(off_div[14]), 
        .B(\un1_sum_adj[14] ), .Y(ADD_32x32_fast_I304_Y_0));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I298_Y_0 (.A(off_div[8]), .B(
        \un1_sum_adj[8] ), .Y(ADD_32x32_fast_I298_Y_0));
    XA1 \off_div_RNO[9]  (.A(N799), .B(ADD_32x32_fast_I299_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[9] ));
    NOR3B \off_div_RNIM95E5[31]  (.A(next_off_div_2_sqmuxa_9), .B(
        next_off_div_2_sqmuxa_8), .C(next_off_div37), .Y(
        next_off_div_2_sqmuxa_11));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y_1 (.A(N622), .B(N637), 
        .C(ADD_32x32_fast_I264_Y_0), .Y(ADD_32x32_fast_I264_Y_1));
    GND GND_i (.Y(GND));
    AND3 un13_nsum_adj_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E[4] ));
    DFN1E1C0 \sum_adj[14]  (.D(\nsum_adj_11[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[14]_net_1 ));
    NOR2 \off_div_RNI6RL4[23]  (.A(off_div[23]), .B(off_div[29]), .Y(
        un1_off_divlto31_9));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I138_Y (.A(N526), .B(N523), 
        .C(N522), .Y(N587));
    OR2 \off_div_RNITECO[4]  (.A(off_div[4]), .B(off_div[3]), .Y(
        un5lto4));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y (.A(
        ADD_32x32_fast_I259_un1_Y_0), .B(N784), .C(
        ADD_32x32_fast_I259_Y_3), .Y(N751));
    OR2 \off_div_RNIVHJ4[13]  (.A(off_div[14]), .B(off_div[13]), .Y(
        un5lto14_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I43_Y (.A(off_div[25]), .B(
        off_div[24]), .C(sum_0_0), .Y(N489));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I123_Y (.A(N507), .B(N511), 
        .Y(N572));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I175_Y (.A(N564), .B(N572), 
        .Y(N630));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I106_Y (.A(N494), .B(N490), 
        .Y(N555));
    MX2 \sum_adj_RNO[10]  (.A(sum_10), .B(I_28_1), .S(sum_1_0), .Y(
        \nsum_adj_11[10] ));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I317_Y (.A(I262_un1_Y), .B(
        ADD_32x32_fast_I262_Y_1), .C(ADD_32x32_fast_I317_Y_0), .Y(
        \un1_off_div_1[27] ));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I11_G0N (.A(sum_1_0), .B(
        \sum_adj[19]_net_1 ), .C(off_div[11]), .Y(N416));
    NOR3C \off_div_RNICHUD1[23]  (.A(un1_off_divlto31_10), .B(
        un1_off_divlto31_9), .C(un1_off_divlt31), .Y(
        un1_off_divlto31_20));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I314_Y_0 (.A(off_div[24]), 
        .B(sum_39), .Y(ADD_32x32_fast_I314_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I271_un1_Y_0 (.A(N586), .B(
        N594), .C(N601), .Y(ADD_32x32_fast_I271_un1_Y_0));
    DFN1E0C0 \off_div[21]  (.D(\next_off_div[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[21]));
    XA1 \off_div_RNO[11]  (.A(N793), .B(ADD_32x32_fast_I301_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[11] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I42_Y (.A(off_div[25]), .B(
        off_div[24]), .C(sum_0_0), .Y(N488));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y (.A(
        ADD_32x32_fast_I263_un1_Y_0), .B(N796), .C(
        ADD_32x32_fast_I263_Y_1), .Y(N759));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I248_Y (.A(N654), .B(N538), 
        .C(N653), .Y(N799));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I301_Y_0 (.A(sum_1_0), .B(
        \sum_adj[19]_net_1 ), .C(off_div[11]), .Y(
        ADD_32x32_fast_I301_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y (.A(
        ADD_32x32_fast_I260_un1_Y_0), .B(N787), .C(
        ADD_32x32_fast_I260_Y_2), .Y(N753));
    AND3 un13_nsum_adj_I_68 (.A(\DWACT_FINC_E[34] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[29] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I306_Y_0 (.A(off_div[16]), 
        .B(sum_39), .Y(ADD_32x32_fast_I306_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I155_Y_0 (.A(off_div[29]), .B(
        off_div[30]), .C(sum_0_0), .Y(ADD_32x32_fast_I155_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I80_Y (.A(N398), .B(N402), .C(
        N401), .Y(N526));
    DFN1E1C0 \sum_adj[13]  (.D(\nsum_adj_11[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[13]_net_1 ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I265_un1_Y_0 (.A(N624), .B(
        N640), .Y(ADD_32x32_fast_I265_un1_Y_0));
    NOR2A \state_RNIVSHN[0]  (.A(state[1]), .B(state[0]), .Y(
        \state_d_0[2] ));
    NOR3A \off_div_RNIMR69[11]  (.A(un1_off_divlto31_2), .B(
        off_div[10]), .C(off_div[11]), .Y(un1_off_divlto31_12));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I170_Y (.A(N567), .B(N560), 
        .C(N559), .Y(N625));
    DFN1E0C0 \off_div[5]  (.D(\next_off_div[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[5]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I7_G0N (.A(\un1_sum_adj[7] )
        , .B(off_div[7]), .Y(N404));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I57_Y (.A(off_div[17]), .B(
        off_div[18]), .C(sum_1_0), .Y(N503));
    XOR2 \state_RNO[1]  (.A(state[1]), .B(state[0]), .Y(N_311_i));
    NOR3A \off_div_RNITB4J1[26]  (.A(un1_off_divlto31_0), .B(
        off_div[26]), .C(un5lto9), .Y(un1_off_divlto31_17));
    NOR3 un13_nsum_adj_I_18 (.A(sum_4), .B(sum_3), .C(sum_5), .Y(
        \DWACT_FINC_E[2] ));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I308_Y (.A(I236_un1_Y), .B(
        ADD_32x32_fast_I271_Y_0), .C(ADD_32x32_fast_I308_Y_0), .Y(
        \un1_off_div_1[18] ));
    MX2 \sum_adj_RNO[11]  (.A(sum_11), .B(I_32_1), .S(sum_1_0), .Y(
        \nsum_adj_11[11] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I321_Y_0 (.A(off_div[31]), 
        .B(sum_39), .Y(ADD_32x32_fast_I321_Y_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I116_Y (.A(N500), .B(N504), 
        .Y(N565));
    NOR2 un13_nsum_adj_I_38 (.A(sum_12), .B(sum_13), .Y(
        \DWACT_FINC_E[8] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I311_Y_0 (.A(off_div[21]), 
        .B(sum_39), .Y(ADD_32x32_fast_I311_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I269_Y_0 (.A(N647), .B(N632), 
        .C(N631), .Y(ADD_32x32_fast_I269_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I81_Y (.A(off_div[5]), .B(
        \un1_sum_adj[5] ), .C(N402), .Y(N527));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I245_Y (.A(N648), .B(N663), 
        .C(N647), .Y(N790));
    MX2 \sum_adj_RNO[12]  (.A(sum_12), .B(I_35_1), .S(sum_1_0), .Y(
        \nsum_adj_11[12] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I316_Y_0 (.A(off_div[26]), 
        .B(sum_39), .Y(ADD_32x32_fast_I316_Y_0));
    XNOR2 un13_nsum_adj_I_46 (.A(sum_16), .B(N_9), .Y(I_46_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I70_Y (.A(N413), .B(N417), .C(
        N416), .Y(N516));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I192_Y (.A(N589), .B(N582), 
        .C(N581), .Y(N647));
    XNOR2 un13_nsum_adj_I_28 (.A(sum_10), .B(N_15), .Y(I_28_1));
    DFN1E0C0 \off_div[30]  (.D(\next_off_div[30] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[30]));
    NOR2 \off_div_RNI1KJ4[14]  (.A(off_div[15]), .B(off_div[14]), .Y(
        un1_off_divlto31_4));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I129_Y (.A(N513), .B(N517), 
        .Y(N578));
    NOR3A \off_div_RNI6C79[16]  (.A(un1_off_divlto31_4), .B(
        off_div[17]), .C(off_div[16]), .Y(un1_off_divlto31_13));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I182_Y (.A(N579), .B(N572), 
        .C(N571), .Y(N637));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I127_Y (.A(N515), .B(N511), 
        .Y(N576));
    VCC VCC_i (.Y(VCC));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I249_Y (.A(I249_un1_Y), .B(
        N655), .Y(N802));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I0_G0N (.A(off_div[0]), .B(
        sum_39), .Y(N383));
    AO1C \state_RNI3P9DA[1]  (.A(un5lt31), .B(next_off_div_2_sqmuxa_11)
        , .C(state[1]), .Y(un1_state_2));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I196_un1_Y (.A(N593), .B(
        N586), .Y(I196_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I45_Y (.A(off_div[23]), .B(
        off_div[24]), .C(sum_0_0), .Y(N491));
    AND3 un13_nsum_adj_I_52 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[12] ), .Y(N_7));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I111_Y (.A(N495), .B(N499), 
        .Y(N560));
    NOR2 \off_div_RNI9SJ4[18]  (.A(off_div[19]), .B(off_div[18]), .Y(
        un1_off_divlto31_6));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I71_Y (.A(off_div[10]), .B(
        \un1_sum_adj[10] ), .C(N417), .Y(N517));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I9_G0N (.A(sum_2_0), .B(
        \sum_adj[17]_net_1 ), .C(off_div[9]), .Y(N410));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I228_un1_Y (.A(N643), .B(
        N628), .Y(I228_un1_Y));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I307_Y_0 (.A(off_div[17]), 
        .B(sum_39), .Y(ADD_32x32_fast_I307_Y_0));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I2_G0N (.A(sum_2_0), .B(
        \sum_adj[10]_net_1 ), .C(off_div[2]), .Y(N389));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I148_Y (.A(N536), .B(N533), 
        .C(N532), .Y(N597));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I48_Y (.A(off_div[21]), .B(
        off_div[22]), .C(sum_0_0), .Y(N494));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I260_un1_Y_0 (.A(N614), .B(
        N630), .Y(ADD_32x32_fast_I260_un1_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I268_un1_Y (.A(N630), .B(
        N646), .C(N661), .Y(I268_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_3 (.A(N612), .B(N627), 
        .C(ADD_32x32_fast_I259_Y_2), .Y(ADD_32x32_fast_I259_Y_3));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I266_un1_Y_0 (.A(N642), .B(
        N626), .Y(ADD_32x32_fast_I266_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I67_Y (.A(N423), .B(N420), 
        .Y(N513));
    XNOR2 un13_nsum_adj_I_70 (.A(sum_23), .B(N_2), .Y(I_70_1));
    NOR3C \off_div_RNIG8K02[20]  (.A(un1_off_divlto31_15), .B(
        un1_off_divlto31_14), .C(un1_off_divlto31_20), .Y(
        un1_off_divlto31_22));
    NOR3A un13_nsum_adj_I_66 (.A(\DWACT_FINC_E[15] ), .B(sum_21), .C(
        sum_22), .Y(\DWACT_FINC_E[33] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I193_Y (.A(N590), .B(N582), 
        .Y(N648));
    NOR2 \off_div_RNI9UL4[27]  (.A(off_div[28]), .B(off_div[27]), .Y(
        un1_off_divlto31_10));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I5_G0N (.A(\un1_sum_adj[5] )
        , .B(off_div[5]), .Y(N398));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I317_Y_0 (.A(off_div[27]), 
        .B(sum_39), .Y(ADD_32x32_fast_I317_Y_0));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y_1 (.A(N486), .B(N482), 
        .C(N555), .Y(ADD_32x32_fast_I260_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I243_Y (.A(N644), .B(N659), 
        .C(N643), .Y(N784));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I296_Y_0 (.A(sum_0_0), .B(
        \sum_adj[14]_net_1 ), .C(off_div[6]), .Y(
        ADD_32x32_fast_I296_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I183_Y (.A(N580), .B(N572), 
        .Y(N638));
    MX2 \sum_adj_RNO[8]  (.A(sum_8), .B(I_23_5), .S(sum_2_0), .Y(
        \nsum_adj_11[8] ));
    XA1 \off_div_RNO[6]  (.A(N659), .B(ADD_32x32_fast_I296_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[6] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I124_Y (.A(N512), .B(N509), 
        .C(N508), .Y(N573));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I273_Y_0 (.A(
        ADD_32x32_fast_I273_un1_Y_0), .B(N640), .C(N639), .Y(
        ADD_32x32_fast_I273_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I157_Y_0 (.A(off_div[28]), .B(
        off_div[29]), .C(sum_2_0), .Y(ADD_32x32_fast_I157_Y_0));
    OA1 \off_div_RNIKEI41[1]  (.A(off_div[1]), .B(off_div[0]), .C(
        off_div[2]), .Y(un5lt4));
    NOR3B un13_nsum_adj_I_36 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .C(sum_12), .Y(N_12));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I242_Y (.A(N642), .B(N657), 
        .C(N641), .Y(N781));
    DFN1E0C0 \off_div[1]  (.D(\next_off_div[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[1]));
    NOR2 un13_nsum_adj_I_47 (.A(sum_15), .B(sum_16), .Y(
        \DWACT_FINC_E[11] ));
    XA1 \off_div_RNO[8]  (.A(N802), .B(ADD_32x32_fast_I298_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[8] ));
    NOR3C \state_RNINJ405[0]  (.A(state[1]), .B(state[0]), .C(
        next_off_div37), .Y(next_off_div_0_sqmuxa));
    XNOR2 un13_nsum_adj_I_26 (.A(sum_9), .B(N_16), .Y(I_26_1));
    OR3 \off_div_RNIQV69[11]  (.A(off_div[12]), .B(off_div[11]), .C(
        un5lto14_1), .Y(un5lto14_2));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I102_Y (.A(N486), .B(N490), 
        .Y(N551));
    XNOR2 un13_nsum_adj_I_43 (.A(sum_15), .B(N_10), .Y(I_43_1));
    XOR2 \sum_adj_RNI4FFU[16]  (.A(\sum_adj[16]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[8] ));
    MX2 \off_div_RNO[19]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[19] ), .S(\state_d[2] ), .Y(\next_off_div[19] ));
    DFN1E0C0 \off_div[10]  (.D(\next_off_div[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[10]));
    MX2 \off_div_RNO[10]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[10] ), .S(\state_d[2] ), .Y(\next_off_div[10] ));
    XOR2 \sum_adj_RNI3EFU[15]  (.A(\sum_adj[15]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[7] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I125_Y (.A(N509), .B(N513), 
        .Y(N574));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y_0 (.A(N553), .B(N561), 
        .Y(ADD_32x32_fast_I263_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I178_Y (.A(N575), .B(N568), 
        .C(N567), .Y(N633));
    NOR3C \off_div_RNIPJI52[11]  (.A(un1_off_divlto31_13), .B(
        un1_off_divlto31_12), .C(un1_off_divlto31_17), .Y(
        un1_off_divlto31_21));
    DFN1E1C0 \sum_adj[12]  (.D(\nsum_adj_11[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[12]_net_1 ));
    NOR3 un13_nsum_adj_I_50 (.A(sum_16), .B(sum_15), .C(sum_17), .Y(
        \DWACT_FINC_E[12] ));
    MX2 \sum_adj_RNO[17]  (.A(sum_17), .B(I_49_1), .S(sum_1_0), .Y(
        \nsum_adj_11[17] ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I297_Y (.A(\un1_sum_adj[7] ), 
        .B(off_div[7]), .C(N657), .Y(\un1_off_div_1[7] ));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I269_un1_Y (.A(N632), .B(
        N648), .C(N663), .Y(I269_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I136_Y (.A(N524), .B(N521), 
        .C(N520), .Y(N585));
    XA1 \off_div_RNO[16]  (.A(N779), .B(ADD_32x32_fast_I306_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[16] ));
    MX2 \off_div_RNO[0]  (.A(next_off_div_0_sqmuxa), .B(
        \un1_off_div_1[0] ), .S(\state_d_0[2] ), .Y(\next_off_div[0] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I199_Y (.A(N596), .B(N588), 
        .Y(N654));
    NOR3B \state_RNINJ405_0[0]  (.A(state[1]), .B(state[0]), .C(
        next_off_div37), .Y(next_off_div_1_sqmuxa));
    XA1 \off_div_RNO[23]  (.A(N765), .B(ADD_32x32_fast_I313_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[23] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I264_un1_Y_0 (.A(N622), .B(
        N638), .Y(ADD_32x32_fast_I264_un1_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I87_Y (.A(off_div[3]), .B(
        \un1_sum_adj[3] ), .C(N390), .Y(N533));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I189_Y (.A(N586), .B(N578), 
        .Y(N644));
    MX2 \off_div_RNO[18]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[18] ), .S(\state_d[2] ), .Y(\next_off_div[18] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I38_Y (.A(off_div[26]), .B(
        off_div[27]), .C(sum_0_0), .Y(N484));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I187_Y (.A(N584), .B(N576), 
        .Y(N642));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I273_Y (.A(N655), .B(N640), 
        .C(ADD_32x32_fast_I273_Y_0), .Y(N779));
    NOR3 un13_nsum_adj_I_67 (.A(sum_1_d0), .B(sum_0_d0), .C(sum_2_d0), 
        .Y(\DWACT_FINC_E[34] ));
    XA1 \off_div_RNO[25]  (.A(N761), .B(ADD_32x32_fast_I315_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[25] ));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I112_Y (.A(N500), .B(N496), 
        .Y(N561));
    XOR2 \sum_adj_RNIV9FU[11]  (.A(\sum_adj[11]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[3] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I14_G0N (.A(
        \un1_sum_adj[14] ), .B(off_div[14]), .Y(N425));
    DFN1E0C0 \off_div[12]  (.D(\next_off_div[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[12]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I271_Y_0 (.A(
        ADD_32x32_fast_I271_un1_Y_0), .B(N636), .C(N635), .Y(
        ADD_32x32_fast_I271_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I161_Y (.A(N485), .B(N489), 
        .C(N558), .Y(N616));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I103_Y (.A(N487), .B(N491), 
        .Y(N552));
    DFN1E0C0 \off_div[0]  (.D(\next_off_div[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[0]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I131_Y (.A(N519), .B(N515), 
        .Y(N580));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I120_Y (.A(N508), .B(N505), 
        .C(N504), .Y(N569));
    NOR2A un13_nsum_adj_I_63 (.A(\DWACT_FINC_E[15] ), .B(sum_21), .Y(
        \DWACT_FINC_E[16] ));
    OA1 \off_div_RNIDGBJ4[16]  (.A(off_div[16]), .B(un5lt16), .C(
        un5lto20_2), .Y(un5lt31));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I46_Y (.A(off_div[22]), .B(
        off_div[23]), .C(sum_0_0), .Y(N492));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I300_Y_0 (.A(off_div[10]), 
        .B(\un1_sum_adj[10] ), .Y(ADD_32x32_fast_I300_Y_0));
    NOR2A \state_RNIVSHN_0[0]  (.A(state[1]), .B(state[0]), .Y(
        \state_d[2] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I77_Y (.A(off_div[7]), .B(
        \un1_sum_adj[7] ), .C(N408), .Y(N523));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I44_Y (.A(off_div[23]), .B(
        off_div[24]), .C(sum_0_0), .Y(N490));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y_2 (.A(N614), .B(N629), 
        .C(ADD_32x32_fast_I260_Y_1), .Y(ADD_32x32_fast_I260_Y_2));
    DFN1E1C0 \sum_adj[20]  (.D(\nsum_adj_11[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[20]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I53_Y (.A(off_div[20]), .B(
        off_div[19]), .C(sum_1_0), .Y(N499));
    MX2 \off_div_RNO[5]  (.A(next_off_div_0_sqmuxa), .B(
        \un1_off_div_1[5] ), .S(\state_d_0[2] ), .Y(\next_off_div[5] ));
    XNOR2 un13_nsum_adj_I_37 (.A(sum_13), .B(N_12), .Y(I_37_1));
    XA1 \off_div_RNO[2]  (.A(N601), .B(ADD_32x32_fast_I292_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[2] ));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I6_G0N (.A(sum_2_0), .B(
        \sum_adj[14]_net_1 ), .C(off_div[6]), .Y(N401));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I247_un1_Y (.A(N586), .B(
        N594), .C(N601), .Y(I247_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I151_Y (.A(N537), .B(
        \un1_sum_adj[0] ), .C(N536), .Y(N601));
    DFN1E0C0 \off_div[6]  (.D(\next_off_div[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[6]));
    NOR3 un13_nsum_adj_I_33 (.A(sum_10), .B(sum_9), .C(sum_11), .Y(
        \DWACT_FINC_E[7] ));
    DFN1E1C0 \sum_adj[17]  (.D(\nsum_adj_11[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[17]_net_1 ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I320_Y_0 (.A(off_div[30]), 
        .B(sum_39), .Y(ADD_32x32_fast_I320_Y_0));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I305_Y (.A(\un1_sum_adj[15] )
        , .B(off_div[15]), .C(N781), .Y(\un1_off_div_1[15] ));
    NOR3A un13_nsum_adj_I_27 (.A(\DWACT_FINC_E[4] ), .B(sum_8), .C(
        sum_9), .Y(N_15));
    NOR2 \off_div_RNI3LCO[6]  (.A(off_div[6]), .B(off_div[7]), .Y(
        un1_off_divlto31_0));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I310_Y_0 (.A(off_div[20]), 
        .B(sum_39), .Y(ADD_32x32_fast_I310_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I270_Y_0 (.A(N649), .B(N634), 
        .C(N633), .Y(ADD_32x32_fast_I270_Y_0));
    NOR2B \off_div_RNIDOC9[30]  (.A(un1_off_divlto31_10), .B(
        next_off_div_2_sqmuxa_5), .Y(next_off_div_2_sqmuxa_8));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I230_un1_Y (.A(N645), .B(
        N630), .Y(I230_un1_Y));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I52_Y (.A(off_div[19]), .B(
        off_div[20]), .C(sum_0_0), .Y(N498));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I204_Y (.A(I204_un1_Y), .B(
        N595), .Y(N661));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I263_un1_Y_0 (.A(N620), .B(
        N636), .Y(ADD_32x32_fast_I263_un1_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I194_Y (.A(N591), .B(N584), 
        .C(N583), .Y(N649));
    XNOR2 un13_nsum_adj_I_23 (.A(sum_8), .B(N_17), .Y(I_23_5));
    XNOR2 un13_nsum_adj_I_59 (.A(sum_20), .B(N_5), .Y(I_59_1));
    DFN1E0C0 \off_div[20]  (.D(\next_off_div[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[20]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I113_Y (.A(N501), .B(N497), 
        .Y(N562));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I184_Y (.A(I184_un1_Y), .B(
        N573), .Y(N639));
    NOR3 un13_nsum_adj_I_41 (.A(sum_13), .B(sum_12), .C(sum_14), .Y(
        \DWACT_FINC_E[9] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_0 (.A(off_div[29]), .B(
        off_div[28]), .C(sum_1_0), .Y(ADD_32x32_fast_I259_Y_0));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I294_Y_0 (.A(sum_2_0), .B(
        \sum_adj[12]_net_1 ), .C(off_div[4]), .Y(
        ADD_32x32_fast_I294_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I236_un1_Y (.A(N651), .B(
        N636), .Y(I236_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I10_G0N (.A(
        \un1_sum_adj[10] ), .B(off_div[10]), .Y(N413));
    XA1 \off_div_RNO[21]  (.A(N769), .B(ADD_32x32_fast_I311_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[21] ));
    NOR2 \off_div_RNI0LL4[22]  (.A(off_div[24]), .B(off_div[22]), .Y(
        un1_off_divlto31_8));
    DFN1E0C0 \off_div[18]  (.D(\next_off_div[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[18]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I262_un1_Y_0 (.A(N618), .B(
        N634), .Y(ADD_32x32_fast_I262_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I109_Y (.A(N497), .B(N493), 
        .Y(N558));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I146_Y (.A(N534), .B(N531), 
        .C(N530), .Y(N595));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I107_Y (.A(N495), .B(N491), 
        .Y(N556));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I195_Y (.A(N592), .B(N584), 
        .Y(N650));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I63_Y (.A(N426), .B(N429), 
        .Y(N509));
    NOR3B un13_nsum_adj_I_55 (.A(\DWACT_FINC_E[13] ), .B(
        \DWACT_FINC_E[28] ), .C(sum_18), .Y(N_6));
    DFN1E0C0 \off_div[22]  (.D(\next_off_div[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[22]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I185_Y (.A(N582), .B(N574), 
        .Y(N640));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I90_Y (.A(N383), .B(N387), .C(
        N386), .Y(N536));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I55_Y (.A(off_div[19]), .B(
        off_div[18]), .C(sum_1_0), .Y(N501));
    XOR2 \sum_adj_RNI1CFU[13]  (.A(\sum_adj[13]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[5] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I49_Y (.A(off_div[22]), .B(
        off_div[21]), .C(sum_0_0), .Y(N495));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_2 (.A(N484), .B(
        ADD_32x32_fast_I259_Y_0), .C(N553), .Y(ADD_32x32_fast_I259_Y_2)
        );
    XA1 \off_div_RNO[12]  (.A(N790), .B(ADD_32x32_fast_I302_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[12] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I62_Y (.A(N425), .B(N429), .C(
        N428), .Y(N508));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y (.A(
        ADD_32x32_fast_I261_un1_Y_0), .B(N790), .C(
        ADD_32x32_fast_I261_Y_2), .Y(N755));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I141_Y (.A(N525), .B(N529), 
        .Y(N590));
    AND3 un13_nsum_adj_I_61 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[15] ), .Y(N_4));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I36_Y (.A(off_div[27]), .B(
        off_div[28]), .C(sum_0_0), .Y(N482));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I58_Y (.A(off_div[17]), .B(
        off_div[16]), .C(sum_1_0), .Y(N504));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I292_Y_0 (.A(sum_0_0), .B(
        \sum_adj[10]_net_1 ), .C(off_div[2]), .Y(
        ADD_32x32_fast_I292_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I91_Y (.A(sum_2_0), .B(
        off_div[0]), .C(N387), .Y(N537));
    DFN1E0C0 \off_div[17]  (.D(\next_off_div[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[17]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I119_Y (.A(N503), .B(N507), 
        .Y(N568));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I190_Y (.A(N587), .B(N580), 
        .C(N579), .Y(N645));
    AND3 un13_nsum_adj_I_54 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[9] ), .C(\DWACT_FINC_E[12] ), .Y(
        \DWACT_FINC_E[13] ));
    MX2 \sum_adj_RNO[23]  (.A(sum_23), .B(I_70_1), .S(sum_2_0), .Y(
        \nsum_adj_11[23] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I117_Y (.A(N501), .B(N505), 
        .Y(N566));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I132_Y (.A(N520), .B(N517), 
        .C(N516), .Y(N581));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I180_Y (.A(N577), .B(N570), 
        .C(N569), .Y(N635));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I128_Y (.A(N516), .B(N513), 
        .C(N512), .Y(N577));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I104_Y (.A(N492), .B(N488), 
        .Y(N553));
    NOR3A un13_nsum_adj_I_31 (.A(\DWACT_FINC_E[6] ), .B(sum_9), .C(
        sum_10), .Y(N_14));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I9_P0N (.A(sum_2_0), .B(
        \sum_adj[17]_net_1 ), .C(off_div[9]), .Y(N411));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I15_G0N (.A(
        \un1_sum_adj[15] ), .B(off_div[15]), .Y(N428));
    NOR2 \off_div_RNI4QM4[30]  (.A(off_div[30]), .B(off_div[29]), .Y(
        next_off_div_2_sqmuxa_5));
    NOR2 un13_nsum_adj_I_21 (.A(sum_6), .B(sum_7), .Y(
        \DWACT_FINC_E[3] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I295_Y_0 (.A(off_div[5]), .B(
        \un1_sum_adj[5] ), .Y(ADD_32x32_fast_I295_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I176_Y (.A(N573), .B(N566), 
        .C(N565), .Y(N631));
    DFN1E0C0 \off_div[28]  (.D(\next_off_div[28] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[28]));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I83_Y (.A(off_div[5]), .B(
        \un1_sum_adj[5] ), .C(N396), .Y(N529));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I65_Y (.A(N423), .B(N426), 
        .Y(N511));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I246_un1_Y (.A(N650), .B(
        N599), .Y(I246_un1_Y));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I12_P0N (.A(\un1_sum_adj[12] )
        , .B(off_div[12]), .Y(N420));
    DFN1C0 \state[1]  (.D(N_311_i), .CLK(clk_c), .CLR(n_rst_c), .Q(
        state[1]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I15_P0N (.A(\un1_sum_adj[15] )
        , .B(off_div[15]), .Y(N429));
    XA1 \off_div_RNO[31]  (.A(N749), .B(ADD_32x32_fast_I321_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[31] ));
    XA1 \off_div_RNO[14]  (.A(N784), .B(ADD_32x32_fast_I304_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[14] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I105_Y (.A(N493), .B(N489), 
        .Y(N554));
    AND3 un13_nsum_adj_I_42 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[9] ), .Y(N_10));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I163_Y (.A(N560), .B(N552), 
        .Y(N618));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I133_Y (.A(N517), .B(N521), 
        .Y(N582));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I68_Y (.A(N416), .B(N420), .C(
        N419), .Y(N514));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I114_Y (.A(N502), .B(N498), 
        .Y(N563));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I261_un1_Y_0 (.A(N616), .B(
        N632), .Y(ADD_32x32_fast_I261_un1_Y_0));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I82_Y (.A(N395), .B(
        off_div[5]), .C(\un1_sum_adj[5] ), .Y(N528));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I171_Y (.A(N560), .B(N568), 
        .Y(N626));
    MX2 \sum_adj_RNO[14]  (.A(sum_14), .B(I_40_1), .S(sum_1_0), .Y(
        \nsum_adj_11[14] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I40_Y (.A(off_div[26]), .B(
        off_div[25]), .C(sum_0_0), .Y(N486));
    DFN1E1C0 \sum_adj[8]  (.D(\nsum_adj_11[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[8]_net_1 ));
    OR2B \off_div_RNITNI41[5]  (.A(un5lto4), .B(off_div[5]), .Y(
        un1_off_divlt31));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I204_un1_Y (.A(N596), .B(
        N538), .Y(I204_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I12_G0N (.A(
        \un1_sum_adj[12] ), .B(off_div[12]), .Y(N419));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I11_P0N (.A(sum_1_0), .B(
        \sum_adj[19]_net_1 ), .C(off_div[11]), .Y(N417));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I73_Y (.A(off_div[10]), .B(
        \un1_sum_adj[10] ), .C(N411), .Y(N519));
    NOR3A \off_div_RNI6GB9[23]  (.A(next_off_div_2_sqmuxa_3), .B(
        off_div[23]), .C(off_div[24]), .Y(next_off_div_2_sqmuxa_7));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I266_Y_0 (.A(N641), .B(N626), 
        .C(N625), .Y(ADD_32x32_fast_I266_Y_0));
    AND3 un13_nsum_adj_I_58 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[14] ), .Y(N_5));
    OA1B \state_RNO[0]  (.A(state[1]), .B(pwm_enable), .C(state[0]), 
        .Y(\state_ns[0] ));
    DFN1E0C0 \off_div[2]  (.D(\next_off_div[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[2]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I39_Y (.A(off_div[27]), .B(
        off_div[26]), .C(sum_0_0), .Y(N485));
    DFN1E0C0 \off_div[27]  (.D(\next_off_div[27] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[27]));
    MX2 \sum_adj_RNO[18]  (.A(sum_18), .B(I_53_1), .S(sum_1_0), .Y(
        \nsum_adj_11[18] ));
    DFN1E1C0 \sum_adj[15]  (.D(\nsum_adj_11[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[15]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I41_Y (.A(off_div[25]), .B(
        off_div[26]), .C(sum_0_0), .Y(N487));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y (.A(
        ADD_32x32_fast_I264_un1_Y_0), .B(N799), .C(
        ADD_32x32_fast_I264_Y_1), .Y(N761));
    NOR3A \off_div_RNI0BC9[30]  (.A(un1_off_divlto31_8), .B(
        off_div[25]), .C(off_div[30]), .Y(un1_off_divlto31_15));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I72_Y (.A(N410), .B(
        off_div[10]), .C(\un1_sum_adj[10] ), .Y(N518));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I295_Y (.A(
        ADD_32x32_fast_I295_Y_0), .B(N661), .Y(\un1_off_div_1[5] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I262_un1_Y (.A(
        ADD_32x32_fast_I262_un1_Y_0), .B(N793), .Y(I262_un1_Y));
    XA1 \off_div_RNO[29]  (.A(N753), .B(ADD_32x32_fast_I319_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[29] ));
    DFN1E0C0 \off_div[14]  (.D(\next_off_div[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[14]));
    DFN1E1C0 \sum_adj[10]  (.D(\nsum_adj_11[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[10]_net_1 ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I302_Y_0 (.A(off_div[12]), 
        .B(\un1_sum_adj[12] ), .Y(ADD_32x32_fast_I302_Y_0));
    MX2 \off_div_RNO[20]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[20] ), .S(\state_d[2] ), .Y(\next_off_div[20] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I300_Y (.A(
        ADD_32x32_fast_I300_Y_0), .B(N796), .Y(\un1_off_div_1[10] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I115_Y (.A(N503), .B(N499), 
        .Y(N564));
    XOR2 \sum_adj_RNIG2CN[20]  (.A(\sum_adj[20]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[12] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I258_un1_Y_0 (.A(N610), .B(
        N626), .Y(ADD_32x32_fast_I258_un1_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I142_Y (.A(N530), .B(N527), 
        .C(N526), .Y(N591));
    XNOR2 un13_nsum_adj_I_62 (.A(sum_21), .B(N_4), .Y(I_62_1));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I56_Y (.A(off_div[18]), .B(
        off_div[17]), .C(sum_1_0), .Y(N502));
    XA1 \off_div_RNO[26]  (.A(N759), .B(ADD_32x32_fast_I316_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[26] ));
    NOR2 \off_div_RNITHL4[21]  (.A(off_div[22]), .B(off_div[21]), .Y(
        next_off_div_2_sqmuxa_1));
    MX2 \sum_adj_RNO[13]  (.A(sum_13), .B(I_37_1), .S(sum_1_0), .Y(
        \nsum_adj_11[13] ));
    DFN1E1C0 \sum_adj[19]  (.D(\nsum_adj_11[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[19]_net_1 ));
    NOR3A \off_div_RNI4C99[20]  (.A(un1_off_divlto31_6), .B(
        off_div[20]), .C(off_div[21]), .Y(un1_off_divlto31_14));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I267_un1_Y (.A(N628), .B(
        N644), .C(N659), .Y(I267_un1_Y));
    MX2 \off_div_RNO[17]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[17] ), .S(\state_d[2] ), .Y(\next_off_div[17] ));
    NOR3C \off_div_RNIHQ5S[21]  (.A(next_off_div_2_sqmuxa_1), .B(
        next_off_div_2_sqmuxa_0), .C(next_off_div_2_sqmuxa_7), .Y(
        next_off_div_2_sqmuxa_9));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I54_Y (.A(off_div[18]), .B(
        off_div[19]), .C(sum_1_0), .Y(N500));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I267_Y (.A(I228_un1_Y), .B(
        N627), .C(I267_un1_Y), .Y(N767));
    DFN1E0P0 \off_div[4]  (.D(\next_off_div[4] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2), .Q(off_div[4]));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I303_Y_0 (.A(sum_2_0), .B(
        \sum_adj[21]_net_1 ), .C(off_div[13]), .Y(
        ADD_32x32_fast_I303_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I169_Y (.A(N566), .B(N558), 
        .Y(N624));
    DFN1E0C0 \off_div[19]  (.D(\next_off_div[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[19]));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I85_Y (.A(off_div[3]), .B(
        \un1_sum_adj[3] ), .C(N396), .Y(N531));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I312_Y_0 (.A(off_div[22]), 
        .B(sum_39), .Y(ADD_32x32_fast_I312_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I139_Y (.A(N523), .B(N527), 
        .Y(N588));
    XA1 \off_div_RNO[28]  (.A(N755), .B(ADD_32x32_fast_I318_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[28] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I167_Y (.A(N564), .B(N556), 
        .Y(N622));
    NOR2 \off_div_RNI5QL4[25]  (.A(off_div[26]), .B(off_div[25]), .Y(
        next_off_div_2_sqmuxa_3));
    DFN1E0C0 \off_div[16]  (.D(\next_off_div[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[16]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I8_P0N (.A(\un1_sum_adj[8] ), 
        .B(off_div[8]), .Y(N408));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I198_Y (.A(N595), .B(N588), 
        .C(N587), .Y(N653));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I137_Y (.A(N525), .B(N521), 
        .Y(N586));
    DFN1E0P0 \off_div[8]  (.D(\next_off_div[8] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2), .Q(off_div[8]));
    XNOR2 un13_nsum_adj_I_32 (.A(sum_11), .B(N_14), .Y(I_32_1));
    XOR2 \sum_adj_RNIJ5CN[23]  (.A(\sum_adj[23]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[15] ));
    NOR2 \off_div_RNITFJ4[12]  (.A(off_div[12]), .B(off_div[13]), .Y(
        un1_off_divlto31_2));
    XOR2 \sum_adj_RNIN8BN[18]  (.A(\sum_adj[18]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[10] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I188_Y (.A(N585), .B(N578), 
        .C(N577), .Y(N643));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I16_P0N (.A(off_div[16]), .B(
        sum_39), .Y(N432));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I110_Y (.A(N498), .B(N494), 
        .Y(N559));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I88_Y (.A(N386), .B(N390), .C(
        N389), .Y(N534));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0 (.A(off_div[30]), .B(
        off_div[29]), .C(sum_0_0), .Y(ADD_32x32_fast_I258_Y_0));
    AND3 un13_nsum_adj_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_17));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I310_Y (.A(I269_un1_Y), .B(
        ADD_32x32_fast_I269_Y_0), .C(ADD_32x32_fast_I310_Y_0), .Y(
        \un1_off_div_1[20] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y_2 (.A(N616), .B(N631), 
        .C(ADD_32x32_fast_I261_Y_1), .Y(ADD_32x32_fast_I261_Y_2));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I159_Y (.A(N483), .B(N487), 
        .C(N556), .Y(N614));
    XNOR2 un13_nsum_adj_I_40 (.A(sum_14), .B(N_11), .Y(I_40_1));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I313_Y_0 (.A(off_div[23]), 
        .B(sum_39), .Y(ADD_32x32_fast_I313_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I157_Y (.A(N485), .B(
        ADD_32x32_fast_I157_Y_0), .C(N554), .Y(N612));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I75_Y (.A(N411), .B(N408), 
        .Y(N521));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I293_Y (.A(
        ADD_32x32_fast_I293_Y_0), .B(N599), .Y(\un1_off_div_1[3] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I143_Y (.A(N527), .B(N531), 
        .Y(N592));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I259_un1_Y_0 (.A(N612), .B(
        N628), .Y(ADD_32x32_fast_I259_un1_Y_0));
    DFN1E0C0 \off_div[3]  (.D(\next_off_div[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[3]));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I290_Y (.A(sum_0_0), .B(
        off_div[0]), .C(\un1_sum_adj[0] ), .Y(\un1_off_div_1[0] ));
    XNOR2 un13_nsum_adj_I_56 (.A(sum_19), .B(N_6), .Y(I_56_1));
    XOR2 \sum_adj_RNII4CN[22]  (.A(\sum_adj[22]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[14] ));
    MX2 \off_div_RNO[7]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[7] ), .S(\state_d_0[2] ), .Y(\next_off_div[7] ));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I78_Y (.A(N401), .B(
        off_div[7]), .C(\un1_sum_adj[7] ), .Y(N524));
    DFN1E1C0 \sum_adj[21]  (.D(\nsum_adj_11[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[21]_net_1 ));
    NOR3C \off_div_RNI9G89[17]  (.A(off_div[18]), .B(off_div[17]), .C(
        un5lto20_1), .Y(un5lto20_2));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_3 (.A(N610), .B(N625), 
        .C(ADD_32x32_fast_I258_Y_2), .Y(ADD_32x32_fast_I258_Y_3));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I66_Y (.A(N419), .B(N423), .C(
        N422), .Y(N512));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I270_un1_Y (.A(N634), .B(
        N650), .C(N599), .Y(I270_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I8_G0N (.A(\un1_sum_adj[8] )
        , .B(off_div[8]), .Y(N407));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I224_un1_Y (.A(N624), .B(
        N639), .Y(I224_un1_Y));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I299_Y_0 (.A(sum_2_0), .B(
        \sum_adj[17]_net_1 ), .C(off_div[9]), .Y(
        ADD_32x32_fast_I299_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I1_G0N (.A(\un1_sum_adj[1] )
        , .B(off_div[1]), .Y(N386));
    XA1 \off_div_RNO[4]  (.A(N663), .B(ADD_32x32_fast_I294_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[4] ));
    DFN1E0C0 \off_div[24]  (.D(\next_off_div[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[24]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I64_Y (.A(N422), .B(N426), .C(
        N425), .Y(N510));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I205_Y (.A(N598), .B(
        \un1_sum_adj[0] ), .C(N597), .Y(N663));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I172_Y (.A(N569), .B(N562), 
        .C(N561), .Y(N627));
    NOR2A \state_RNIVSHN_1[0]  (.A(state[0]), .B(state[1]), .Y(
        state_176_d));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I3_G0N (.A(\un1_sum_adj[3] )
        , .B(off_div[3]), .Y(N392));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I134_Y (.A(N522), .B(N519), 
        .C(N518), .Y(N583));
    DFN1E1C0 \sum_adj[16]  (.D(\nsum_adj_11[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[16]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I244_Y (.A(N646), .B(N661), 
        .C(N645), .Y(N787));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I238_un1_Y (.A(N653), .B(
        N638), .Y(I238_un1_Y));
    MX2 \sum_adj_RNO[19]  (.A(sum_19), .B(I_56_1), .S(sum_1_0), .Y(
        \nsum_adj_11[19] ));
    XOR2 \sum_adj_RNIMQ5T[9]  (.A(\sum_adj[9]_net_1 ), .B(sum_39), .Y(
        \un1_sum_adj[1] ));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I6_P0N (.A(sum_2_0), .B(
        \sum_adj[14]_net_1 ), .C(off_div[6]), .Y(N402));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y_1 (.A(N484), .B(N488), 
        .C(N557), .Y(ADD_32x32_fast_I261_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I126_Y (.A(N514), .B(N511), 
        .C(N510), .Y(N575));
    NOR3 un13_nsum_adj_I_60 (.A(sum_19), .B(sum_18), .C(sum_20), .Y(
        \DWACT_FINC_E[15] ));
    XA1 \off_div_RNO[30]  (.A(N751), .B(ADD_32x32_fast_I320_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[30] ));
    
endmodule


module integral_calc_13s_4_1(
       avg_old,
       avg_new,
       LED_33_0,
       choose,
       LED_5_0,
       LED_c_0,
       choose_0_0,
       LED_15_0,
       LED_12_0,
       average,
       LED_FB,
       LED_FB_i_0,
       calc_avg,
       avg_done,
       n_rst_c,
       clk_c
    );
input  [11:0] avg_old;
input  [11:0] avg_new;
input  LED_33_0;
input  [2:0] choose;
input  LED_5_0;
output LED_c_0;
input  choose_0_0;
input  LED_15_0;
input  LED_12_0;
output [6:2] average;
output [7:0] LED_FB;
output LED_FB_i_0;
input  calc_avg;
output avg_done;
input  n_rst_c;
input  clk_c;

    wire \state_1[0]_net_1 , \state_RNI3U7Q[0]_net_1 , 
        \state_0[0]_net_1 , N427, N339, N342, N435, N330, N327, N437, 
        N324, \un1_next_int[7] , \un1_next_int[2] , \un1_next_int[4] , 
        \un1_next_int[8] , \un1_next_int[3] , ADD_26x26_fast_I253_Y_0, 
        \integ[23]_net_1 , \state[0]_net_1 , ADD_26x26_fast_I255_Y_0, 
        \integ[25]_net_1 , ADD_26x26_fast_I254_Y_0, \integ[24]_net_1 , 
        ADD_26x26_fast_I206_Y_2, N506, N521, ADD_26x26_fast_I206_Y_1, 
        N398, N402, N459, ADD_26x26_fast_I252_Y_0, \integ[22]_net_1 , 
        ADD_26x26_fast_I205_Y_3, N504, N519, ADD_26x26_fast_I205_Y_2, 
        N400, ADD_26x26_fast_I205_Y_0, N457, ADD_26x26_fast_I204_Y_3, 
        N502, N517, ADD_26x26_fast_I204_Y_2, N406, 
        ADD_26x26_fast_I204_Y_1, ADD_26x26_fast_I204_Y_0, 
        ADD_26x26_fast_I251_Y_0, \integ[21]_net_1 , 
        ADD_26x26_fast_I250_Y_0, \integ[20]_net_1 , 
        ADD_26x26_fast_I249_Y_0, \integ[19]_net_1 , 
        ADD_26x26_fast_I207_Y_2, N508, N523, ADD_26x26_fast_I207_Y_1, 
        N404, N461, ADD_26x26_fast_I248_Y_0, \integ[18]_net_1 , 
        ADD_26x26_fast_I246_Y_0, \integ[16]_net_1 , 
        ADD_26x26_fast_I247_Y_0, \integ[17]_net_1 , 
        ADD_26x26_fast_I243_Y_0, ADD_26x26_fast_I241_Y_0, 
        \state_RNINB1R[0]_net_1 , ADD_26x26_fast_I208_Y_1, 
        ADD_26x26_fast_I208_un1_Y_0, N541, ADD_26x26_fast_I208_Y_0, 
        N463, ADD_26x26_fast_I209_Y_1, ADD_26x26_fast_I209_un1_Y_0, 
        N543, ADD_26x26_fast_I209_Y_0, N465, N458, 
        ADD_26x26_fast_I239_Y_0, \un1_next_int[9] , 
        ADD_26x26_fast_I210_Y_1, ADD_26x26_fast_I210_un1_Y_0, N491, 
        ADD_26x26_fast_I210_Y_0, N467, N460, 
        ADD_26x26_fast_I204_un1_Y_0, N518, ADD_26x26_fast_I205_un1_Y_0, 
        N520, ADD_26x26_fast_I240_Y_0, \inf_abs0_m[10] , 
        \un18_next_int_m[10] , ADD_26x26_fast_I212_Y_0, 
        ADD_26x26_fast_I212_un1_Y_0, ADD_26x26_fast_I213_Y_0, 
        ADD_26x26_fast_I213_un1_Y_0, ADD_26x26_fast_I211_Y_1, 
        ADD_26x26_fast_I211_un1_Y_0, N516, ADD_26x26_fast_I211_Y_0, 
        N469, N462, ADD_26x26_fast_I235_Y_0, \un18_next_int_m[5] , 
        \inf_abs0_m[5] , ADD_26x26_fast_I234_Y_0, N512, N528, N510, 
        N526, N476, N484, N514, N482, N490, \un1_next_int[0] , N480, 
        N488, N442, N478, N486, N493, ADD_26x26_fast_I232_Y_0, 
        ADD_26x26_fast_I231_Y_0, \un18_next_int_m[1] , \inf_abs0_m[1] , 
        \integ[1]_net_1 , ADD_26x26_fast_I127_Y_0, 
        ADD_26x26_fast_I230_Y_0, \integ[0]_net_1 , \state[1]_net_1 , 
        ADD_26x26_fast_I125_Y_1, ADD_26x26_fast_I125_Y_0, N399, 
        \un1_integ[20] , I178_un1_Y, \un1_integ[16] , I186_un1_Y, 
        \un1_integ[17] , I184_un1_Y, N407, N403, I204_un1_Y, N533, 
        I194_un1_Y, \un1_integ[19] , I180_un1_Y, 
        ADD_26x26_fast_I230_Y_0_0, \un1_integ[25] , \un1_integ[21] , 
        I176_un1_Y, \un1_integ[18] , I182_un1_Y, \un1_integ[14] , N640, 
        \un1_integ[15] , \integ[15]_net_1 , N637, N401, I205_un1_Y, 
        N658, \un1_integ[24] , \un1_integ[6] , \un1_next_int[6] , N539, 
        \un1_integ[12] , N646, ADD_26x26_fast_I233_Y, \un1_integ[7] , 
        N537, \un1_integ[13] , N525, I190_un1_Y, \un1_integ[23] , 
        I206_un1_Y, ADD_26x26_fast_I232_Y, \un1_integ[10] , N531, 
        I193_un1_Y, \un1_integ[22] , I207_un1_Y, \un1_integ[11] , N529, 
        I192_un1_Y, \un1_integ[9] , \un1_integ[8] , \un1_integ[5] , 
        ADD_26x26_fast_I234_Y, ADD_26x26_fast_I231_Y, N522, N524, N405, 
        \inf_abs0_m[11] , \un18_next_int_m[11] , N_101, N_46, N_38, 
        N_70, N_54, N_62, N535, N489, N481, I163_un1_Y, N527, N479, 
        N430, N426, N338, N431, N336, N333, N439, N321, I150_un1_Y, 
        N473, N424, N421, N420, N474, N425, N345, N477, N470, N417, 
        N429, N440, N436, N323, N441, N318, N433, N432, N428, N335, 
        N332, I74_un1_Y, N317, I112_un1_Y, N434, N483, N438, N320, 
        N326, N329, N350, N351, N341, N344, I114_un1_Y, N485, 
        I121_un1_Y, \inf_abs0_m[3] , \un18_next_int_m[3] , 
        \inf_abs0_m[7] , \un18_next_int_m[7] , \inf_abs0_m[2] , 
        \un18_next_int_m[2] , \inf_abs0_m[6] , \un18_next_int_m[6] , 
        \inf_abs0_m[9] , \un18_next_int_m[9] , \state_RNO_3[1] , 
        \inf_abs0_m[0] , \un18_next_int_m[0] , I195_un1_Y, I154_un1_Y, 
        N416, N353, N415, N357, N414, N422, N348, N347, N418, N354, 
        N410, N411, I152_un1_Y, N475, N468, N464, N423, N471, N419, 
        N472, N408, N413, N412, N409, \inf_abs0_m[8] , 
        \un18_next_int_m[8] , \inf_abs0_m[4] , \un18_next_int_m[4] , 
        I162_un1_Y, N487, N466, GND, VCC;
    
    AO1 un1_integ_0_0_ADD_26x26_fast_I56_Y (.A(N341), .B(N345), .C(
        N344), .Y(N424));
    NOR2A \state_RNI4FT8[1]  (.A(\state[1]_net_1 ), .B(avg_old[8]), .Y(
        \un18_next_int_m[8] ));
    DFN1C0 \state[0]  (.D(\state_RNI3U7Q[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[0]_net_1 ));
    DFN1E0C0 \integ[13]  (.D(\un1_integ[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(LED_FB[6]));
    DFN1E0C0 \integ[24]  (.D(\un1_integ[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[24]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I112_un1_Y (.A(N434), .B(N431), 
        .Y(I112_un1_Y));
    OA1 un1_integ_0_0_ADD_26x26_fast_I61_Y (.A(LED_FB[0]), .B(
        \un1_next_int[7] ), .C(N336), .Y(N429));
    OR2 un1_integ_0_0_ADD_26x26_fast_I7_P0N (.A(LED_FB[0]), .B(
        \un1_next_int[7] ), .Y(N339));
    NOR2A \state_RNIS6T8[1]  (.A(\state[1]_net_1 ), .B(avg_old[0]), .Y(
        \un18_next_int_m[0] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I248_Y_0 (.A(\integ[18]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I248_Y_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I41_Y (.A(\integ[17]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N409));
    OA1 un1_integ_0_0_ADD_26x26_fast_I204_un1_Y (.A(N533), .B(
        I194_un1_Y), .C(ADD_26x26_fast_I204_un1_Y_0), .Y(I204_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I86_Y (.A(N408), .B(N404), .Y(
        N457));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I125_Y_1 (.A(
        ADD_26x26_fast_I125_Y_0), .B(N399), .Y(ADD_26x26_fast_I125_Y_1)
        );
    AO1 un1_integ_0_0_ADD_26x26_fast_I98_Y (.A(N420), .B(N417), .C(
        N416), .Y(N469));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I176_un1_Y (.A(N510), .B(N525), 
        .Y(I176_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I205_un1_Y_0 (.A(N504), .B(N520)
        , .Y(ADD_26x26_fast_I205_un1_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I150_un1_Y (.A(N481), .B(N474), 
        .Y(I150_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I51_Y (.A(N354), .B(N351), .Y(
        N419));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y (.A(
        ADD_26x26_fast_I230_Y_0), .B(\un1_next_int[0] ), .Y(
        ADD_26x26_fast_I230_Y_0_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I253_Y (.A(I206_un1_Y), .B(
        ADD_26x26_fast_I206_Y_2), .C(ADD_26x26_fast_I253_Y_0), .Y(
        \un1_integ[23] ));
    DFN1E0C0 \integ[21]  (.D(\un1_integ[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[21]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I190_un1_Y (.A(N526), .B(N541), 
        .Y(I190_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I146_Y (.A(N477), .B(N470), .C(
        N469), .Y(N523));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I210_un1_Y_0 (.A(N476), .B(N484)
        , .C(N514), .Y(ADD_26x26_fast_I210_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I142_Y (.A(N473), .B(N466), .C(
        N465), .Y(N519));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I231_Y (.A(
        ADD_26x26_fast_I231_Y_0), .B(N442), .Y(ADD_26x26_fast_I231_Y));
    MX2 \un1_integ_0_0_LED_7[4]  (.A(N_46), .B(N_70), .S(choose[0]), 
        .Y(LED_c_0));
    DFN1E0C0 \integ[15]  (.D(\un1_integ[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[15]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I103_Y (.A(N421), .B(N425), .Y(
        N474));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I125_Y (.A(N407), .B(N403), .C(
        ADD_26x26_fast_I125_Y_1), .Y(N502));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_1 (.A(
        ADD_26x26_fast_I209_un1_Y_0), .B(N543), .C(
        ADD_26x26_fast_I209_Y_0), .Y(ADD_26x26_fast_I209_Y_1));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I97_Y (.A(N415), .B(N419), .Y(
        N468));
    AO1 un1_integ_0_0_ADD_26x26_fast_I94_Y (.A(N416), .B(N413), .C(
        N412), .Y(N465));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I151_Y (.A(N474), .B(N482), .Y(
        N528));
    NOR2A \un1_integ_0_0_LED_4[4]  (.A(LED_FB[4]), .B(choose[2]), .Y(
        N_54));
    OR2 un1_integ_0_0_ADD_26x26_fast_I74_Y (.A(I74_un1_Y), .B(N317), 
        .Y(N442));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I238_Y (.A(\un1_next_int[8] ), 
        .B(LED_FB[1]), .C(N658), .Y(\un1_integ[8] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I121_Y (.A(I121_un1_Y), .B(N440), 
        .Y(N493));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I154_un1_Y (.A(N485), .B(N478), 
        .Y(I154_un1_Y));
    OR3 un1_integ_0_0_ADD_26x26_fast_I5_P0N (.A(\un18_next_int_m[5] ), 
        .B(\inf_abs0_m[5] ), .C(average[5]), .Y(N333));
    NOR2A \un1_integ_0_0_LED_5[4]  (.A(LED_33_0), .B(choose[2]), .Y(
        N_62));
    AX1D un1_integ_0_0_ADD_26x26_fast_I246_Y (.A(I186_un1_Y), .B(
        ADD_26x26_fast_I213_Y_0), .C(ADD_26x26_fast_I246_Y_0), .Y(
        \un1_integ[16] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I252_Y_0 (.A(\integ[22]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I252_Y_0));
    DFN1C0 \state_1[0]  (.D(\state_RNI3U7Q[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_1[0]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I39_Y (.A(\integ[18]_net_1 ), .B(
        \integ[17]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N407));
    OA1B un1_integ_0_0_ADD_26x26_fast_I32_Y (.A(\integ[20]_net_1 ), .B(
        \integ[21]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N400));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I194_un1_Y (.A(N480), .B(N488), 
        .C(N442), .Y(I194_un1_Y));
    AO1B un1_integ_0_0_ADD_26x26_fast_I125_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\integ[24]_net_1 ), .C(\state_0[0]_net_1 ), .Y(
        ADD_26x26_fast_I125_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I100_Y (.A(N422), .B(N419), .C(
        N418), .Y(N471));
    OR2 un1_integ_0_0_ADD_26x26_fast_I12_P0N (.A(LED_FB[5]), .B(
        \state[1]_net_1 ), .Y(N354));
    OA1 un1_integ_0_0_ADD_26x26_fast_I10_G0N (.A(\inf_abs0_m[10] ), .B(
        \un18_next_int_m[10] ), .C(LED_FB[3]), .Y(N347));
    DFN1E0C0 \integ[12]  (.D(\un1_integ[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(LED_FB[5]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I109_Y (.A(N427), .B(N431), .Y(
        N480));
    OA1B un1_integ_0_0_ADD_26x26_fast_I205_Y_0 (.A(\integ[22]_net_1 ), 
        .B(\integ[23]_net_1 ), .C(\state_0[0]_net_1 ), .Y(
        ADD_26x26_fast_I205_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I115_Y (.A(N433), .B(N437), .Y(
        N486));
    OR2 \state_RNI9OH81[1]  (.A(\inf_abs0_m[3] ), .B(
        \un18_next_int_m[3] ), .Y(\un1_next_int[3] ));
    NOR2B \state_RNI0V4O[0]  (.A(avg_new[9]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[9] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I12_G0N (.A(LED_FB[5]), .B(
        \state[1]_net_1 ), .Y(N353));
    OR3 un1_integ_0_0_ADD_26x26_fast_I208_Y_0 (.A(N406), .B(N402), .C(
        N463), .Y(ADD_26x26_fast_I208_Y_0));
    NOR2A \un1_integ_0_0_LED_2[4]  (.A(LED_5_0), .B(choose[2]), .Y(
        N_38));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I111_Y (.A(N433), .B(N429), .Y(
        N482));
    NOR2A \state_RNIDV4A[1]  (.A(\state[1]_net_1 ), .B(avg_old[10]), 
        .Y(\un18_next_int_m[10] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I2_P0N (.A(average[2]), .B(
        \un1_next_int[2] ), .Y(N324));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I250_Y_0 (.A(\integ[20]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I250_Y_0));
    MX2 \un1_integ_0_0_LED_3[4]  (.A(N_101), .B(N_38), .S(choose[1]), 
        .Y(N_46));
    DFN1E0C0 \integ[10]  (.D(\un1_integ[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(LED_FB[3]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I180_un1_Y (.A(N514), .B(N529), 
        .Y(I180_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I162_Y (.A(I162_un1_Y), .B(N487), 
        .Y(N541));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I6_G0N (.A(\un1_next_int[6] ), 
        .B(average[6]), .Y(N335));
    AX1D un1_integ_0_0_ADD_26x26_fast_I249_Y (.A(I180_un1_Y), .B(
        ADD_26x26_fast_I210_Y_1), .C(ADD_26x26_fast_I249_Y_0), .Y(
        \un1_integ[19] ));
    GND GND_i (.Y(GND));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I246_Y_0 (.A(\integ[16]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I246_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I6_P0N (.A(\un1_next_int[6] ), .B(
        average[6]), .Y(N336));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I212_un1_Y_0 (.A(N480), .B(N488)
        , .C(N442), .Y(ADD_26x26_fast_I212_un1_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I1_G0N (.A(\un18_next_int_m[1] ), 
        .B(\inf_abs0_m[1] ), .C(\integ[1]_net_1 ), .Y(N320));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I107_Y (.A(N425), .B(N429), .Y(
        N478));
    OA1B un1_integ_0_0_ADD_26x26_fast_I38_Y (.A(\integ[17]_net_1 ), .B(
        \integ[18]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N406));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I209_un1_Y_0 (.A(N512), .B(N528)
        , .Y(ADD_26x26_fast_I209_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_3 (.A(N504), .B(N519), .C(
        ADD_26x26_fast_I205_Y_2), .Y(ADD_26x26_fast_I205_Y_3));
    AX1D un1_integ_0_0_ADD_26x26_fast_I255_Y (.A(I204_un1_Y), .B(
        ADD_26x26_fast_I204_Y_3), .C(ADD_26x26_fast_I255_Y_0), .Y(
        \un1_integ[25] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I204_Y_0 (.A(\integ[24]_net_1 ), 
        .B(\integ[23]_net_1 ), .C(\state_0[0]_net_1 ), .Y(
        ADD_26x26_fast_I204_Y_0));
    NOR2B \state_1_RNI9DKV[0]  (.A(avg_new[2]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[2] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I243_Y (.A(N525), .B(I190_un1_Y), 
        .C(ADD_26x26_fast_I243_Y_0), .Y(\un1_integ[13] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I231_Y_0 (.A(
        \un18_next_int_m[1] ), .B(\inf_abs0_m[1] ), .C(
        \integ[1]_net_1 ), .Y(ADD_26x26_fast_I231_Y_0));
    NOR2A \state_RNIT7T8[1]  (.A(\state[1]_net_1 ), .B(avg_old[1]), .Y(
        \un18_next_int_m[1] ));
    AND2 un1_integ_0_0_ADD_26x26_fast_I69_Y (.A(N324), .B(N327), .Y(
        N437));
    AO1 un1_integ_0_0_ADD_26x26_fast_I62_Y (.A(N332), .B(N336), .C(
        N335), .Y(N430));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I193_un1_Y (.A(N478), .B(N486), 
        .C(N493), .Y(I193_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I152_un1_Y (.A(N483), .B(N476), 
        .Y(I152_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I7_G0N (.A(\un1_next_int[7] ), 
        .B(LED_FB[0]), .Y(N338));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I49_Y (.A(N354), .B(N357), .Y(
        N417));
    OA1B un1_integ_0_0_ADD_26x26_fast_I42_Y (.A(\integ[15]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_1[0]_net_1 ), .Y(N410));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I145_Y (.A(N468), .B(N476), .Y(
        N522));
    OR3 un1_integ_0_0_ADD_26x26_fast_I10_P0N (.A(\inf_abs0_m[10] ), .B(
        \un18_next_int_m[10] ), .C(LED_FB[3]), .Y(N348));
    OR3 un1_integ_0_0_ADD_26x26_fast_I1_P0N (.A(\un18_next_int_m[1] ), 
        .B(\inf_abs0_m[1] ), .C(\integ[1]_net_1 ), .Y(N321));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I184_un1_Y (.A(N533), .B(N518), 
        .Y(I184_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I192_un1_Y (.A(N476), .B(N484), 
        .C(N491), .Y(I192_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I141_Y (.A(N464), .B(N472), .Y(
        N518));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I93_Y (.A(N411), .B(N415), .Y(
        N464));
    AO1B un1_integ_0_0_ADD_26x26_fast_I37_Y (.A(\integ[19]_net_1 ), .B(
        \integ[18]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N405));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I0_G0N (.A(\integ[0]_net_1 ), 
        .B(\state[1]_net_1 ), .Y(N317));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I73_Y (.A(N318), .B(N321), .Y(
        N441));
    AND2 un1_integ_0_0_ADD_26x26_fast_I59_Y (.A(N339), .B(N342), .Y(
        N427));
    AO1 un1_integ_0_0_ADD_26x26_fast_I52_Y (.A(N347), .B(N351), .C(
        N350), .Y(N420));
    NOR2A \state_RNO[1]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 ), 
        .Y(\state_RNO_3[1] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I34_Y (.A(\integ[20]_net_1 ), .B(
        \integ[19]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N402));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I236_Y (.A(\un1_next_int[6] ), 
        .B(average[6]), .C(N539), .Y(\un1_integ[6] ));
    NOR2A \state_RNIE05A[1]  (.A(\state[1]_net_1 ), .B(avg_old[11]), 
        .Y(\un18_next_int_m[11] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I150_Y (.A(I150_un1_Y), .B(N473), 
        .Y(N527));
    DFN1C0 \integ[0]  (.D(ADD_26x26_fast_I230_Y_0_0), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\integ[0]_net_1 ));
    NOR2B \state_1_RNIAEKV[0]  (.A(avg_new[3]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[3] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I120_Y (.A(N439), .B(N442), .C(
        N438), .Y(N491));
    AO1 un1_integ_0_0_ADD_26x26_fast_I104_Y (.A(N426), .B(N423), .C(
        N422), .Y(N475));
    NOR2B \state_RNI9BSG[0]  (.A(avg_new[11]), .B(\state[0]_net_1 ), 
        .Y(\inf_abs0_m[11] ));
    VCC VCC_i (.Y(VCC));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I129_Y (.A(N399), .B(N403), .C(
        N460), .Y(N506));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I113_Y (.A(N435), .B(N431), .Y(
        N484));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I241_Y_0 (.A(LED_FB[4]), .B(
        \state_RNINB1R[0]_net_1 ), .Y(ADD_26x26_fast_I241_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I89_Y (.A(N411), .B(N407), .Y(
        N460));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I68_Y (.A(N323), .B(average[3]), 
        .C(\un1_next_int[3] ), .Y(N436));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_0 (.A(N469), .B(N462), .C(
        N461), .Y(ADD_26x26_fast_I211_Y_0));
    NOR2A \state_RNI1CT8[1]  (.A(\state[1]_net_1 ), .B(avg_old[5]), .Y(
        \un18_next_int_m[5] ));
    INV \integ_RNI2448[12]  (.A(LED_FB[5]), .Y(LED_FB_i_0));
    DFN1C0 \integ[4]  (.D(ADD_26x26_fast_I234_Y), .CLK(clk_c), .CLR(
        n_rst_c), .Q(average[4]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I108_Y (.A(N430), .B(N427), .C(
        N426), .Y(N479));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I3_G0N (.A(\un1_next_int[3] ), 
        .B(average[3]), .Y(N326));
    AO13 un1_integ_0_0_ADD_26x26_fast_I48_Y (.A(LED_FB[6]), .B(N353), 
        .C(\state_1[0]_net_1 ), .Y(N416));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I195_un1_Y (.A(N482), .B(N490), 
        .C(\un1_next_int[0] ), .Y(I195_un1_Y));
    NOR2B \state_1_RNIFJKV[0]  (.A(avg_new[8]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[8] ));
    NOR2B \state_1_RNI8CKV[0]  (.A(avg_new[1]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[1] ));
    OR2 \state_RNI3IH81[1]  (.A(\un18_next_int_m[0] ), .B(
        \inf_abs0_m[0] ), .Y(\un1_next_int[0] ));
    DFN1C0 \integ[3]  (.D(ADD_26x26_fast_I233_Y), .CLK(clk_c), .CLR(
        n_rst_c), .Q(average[3]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I252_Y (.A(I207_un1_Y), .B(
        ADD_26x26_fast_I207_Y_2), .C(ADD_26x26_fast_I252_Y_0), .Y(
        \un1_integ[22] ));
    DFN1E0C0 \integ[6]  (.D(\un1_integ[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[6]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_1 (.A(
        ADD_26x26_fast_I210_un1_Y_0), .B(N491), .C(
        ADD_26x26_fast_I210_Y_0), .Y(ADD_26x26_fast_I210_Y_1));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y (.A(N533), .B(I194_un1_Y), 
        .C(ADD_26x26_fast_I239_Y_0), .Y(\un1_integ[9] ));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I58_Y (.A(N338), .B(LED_FB[1]), 
        .C(\un1_next_int[8] ), .Y(N426));
    AND2 un1_integ_0_0_ADD_26x26_fast_I67_Y (.A(N330), .B(N327), .Y(
        N435));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I253_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I253_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I64_Y (.A(N329), .B(N333), .C(
        N332), .Y(N432));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I204_un1_Y_0 (.A(N502), .B(N518)
        , .Y(ADD_26x26_fast_I204_un1_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I127_Y (.A(N401), .B(
        ADD_26x26_fast_I127_Y_0), .C(N458), .Y(N504));
    AO1 un1_integ_0_0_ADD_26x26_fast_I110_Y (.A(N432), .B(N429), .C(
        N428), .Y(N481));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I211_un1_Y_0 (.A(N478), .B(N486)
        , .C(N493), .Y(ADD_26x26_fast_I211_un1_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I90_Y (.A(N412), .B(N408), .Y(
        N461));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I233_Y (.A(\un1_next_int[3] ), 
        .B(average[3]), .C(N491), .Y(ADD_26x26_fast_I233_Y));
    OA1A un1_integ_0_0_ADD_26x26_fast_I47_Y (.A(\state_1[0]_net_1 ), 
        .B(LED_FB[7]), .C(N357), .Y(N415));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I119_Y (.A(N441), .B(N437), .Y(
        N490));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I70_Y (.A(N320), .B(average[2]), 
        .C(\un1_next_int[2] ), .Y(N438));
    NOR2B \state_1_RNIBFKV[0]  (.A(avg_new[4]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[4] ));
    DFN1E0C0 \integ[5]  (.D(\un1_integ[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[5]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I182_un1_Y (.A(N516), .B(N531), 
        .Y(I182_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I161_Y (.A(N486), .B(N493), .C(
        N485), .Y(N539));
    OA1B un1_integ_0_0_ADD_26x26_fast_I44_Y (.A(\integ[15]_net_1 ), .B(
        LED_FB[7]), .C(\state_1[0]_net_1 ), .Y(N412));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I245_Y (.A(\state_0[0]_net_1 ), 
        .B(\integ[15]_net_1 ), .C(N637), .Y(\un1_integ[15] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I95_Y (.A(N413), .B(N417), .Y(
        N466));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I239_Y_0 (.A(LED_FB[2]), .B(
        \un1_next_int[9] ), .Y(ADD_26x26_fast_I239_Y_0));
    DFN1C0 \integ[2]  (.D(ADD_26x26_fast_I232_Y), .CLK(clk_c), .CLR(
        n_rst_c), .Q(average[2]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I135_Y (.A(N466), .B(N458), .Y(
        N512));
    OR2 un1_integ_0_0_ADD_26x26_fast_I88_Y (.A(N410), .B(N406), .Y(
        N459));
    AX1D un1_integ_0_0_ADD_26x26_fast_I247_Y (.A(I184_un1_Y), .B(
        ADD_26x26_fast_I212_Y_0), .C(ADD_26x26_fast_I247_Y_0), .Y(
        \un1_integ[17] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I143_Y (.A(N466), .B(N474), .Y(
        N520));
    NOR2 \state_RNIJSNG[0]  (.A(\state[1]_net_1 ), .B(\state[0]_net_1 )
        , .Y(avg_done));
    OA1 un1_integ_0_0_ADD_26x26_fast_I57_Y (.A(LED_FB[1]), .B(
        \un1_next_int[8] ), .C(N345), .Y(N425));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I186_un1_Y (.A(N535), .B(N520), 
        .Y(I186_un1_Y));
    DFN1E0C0 \integ[23]  (.D(\un1_integ[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[23]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I8_P0N (.A(LED_FB[1]), .B(
        \un1_next_int[8] ), .Y(N342));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_2 (.A(N506), .B(N521), .C(
        ADD_26x26_fast_I206_Y_1), .Y(ADD_26x26_fast_I206_Y_2));
    AO1 un1_integ_0_0_ADD_26x26_fast_I54_Y (.A(N344), .B(N348), .C(
        N347), .Y(N422));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I131_Y (.A(N405), .B(N401), .C(
        N462), .Y(N508));
    AX1D un1_integ_0_0_ADD_26x26_fast_I254_Y (.A(I205_un1_Y), .B(
        ADD_26x26_fast_I205_Y_3), .C(ADD_26x26_fast_I254_Y_0), .Y(
        \un1_integ[24] ));
    DFN1E0C0 \integ[19]  (.D(\un1_integ[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[19]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I117_Y (.A(N439), .B(N435), .Y(
        N488));
    DFN1E0C0 \integ[17]  (.D(\un1_integ[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[17]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I33_Y (.A(\integ[20]_net_1 ), .B(
        \integ[21]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N401));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I255_Y_0 (.A(\integ[25]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I255_Y_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I127_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\integ[22]_net_1 ), .C(\state_1[0]_net_1 ), .Y(
        ADD_26x26_fast_I127_Y_0));
    DFN1E0C0 \integ[14]  (.D(\un1_integ[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(LED_FB[7]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I87_Y (.A(N405), .B(N409), .Y(
        N458));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y_0 (.A(average[2]), .B(
        \un1_next_int[2] ), .Y(ADD_26x26_fast_I232_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I154_Y (.A(I154_un1_Y), .B(N477), 
        .Y(N531));
    OR2 \state_RNIH0I81[1]  (.A(\inf_abs0_m[7] ), .B(
        \un18_next_int_m[7] ), .Y(\un1_next_int[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I11_G0N (.A(
        \state_RNINB1R[0]_net_1 ), .B(LED_FB[4]), .Y(N350));
    MX2 \un1_integ_0_0_LED_1[4]  (.A(LED_12_0), .B(LED_15_0), .S(
        choose_0_0), .Y(N_101));
    AO1 un1_integ_0_0_ADD_26x26_fast_I140_Y (.A(N471), .B(N464), .C(
        N463), .Y(N517));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I149_Y (.A(N480), .B(N472), .Y(
        N526));
    NOR2B \state_1_RNIEIKV[0]  (.A(avg_new[7]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[7] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I158_Y (.A(N489), .B(N482), .C(
        N481), .Y(N535));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I249_Y_0 (.A(\integ[19]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I249_Y_0));
    DFN1E0C0 \integ[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[25]_net_1 ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I247_Y_0 (.A(\integ[17]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I247_Y_0));
    NOR2B \state_RNI8ASG[0]  (.A(avg_new[10]), .B(\state[0]_net_1 ), 
        .Y(\inf_abs0_m[10] ));
    NOR2A \state_RNI0BT8[1]  (.A(\state[1]_net_1 ), .B(avg_old[4]), .Y(
        \un18_next_int_m[4] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y_0 (.A(\integ[0]_net_1 ), 
        .B(\state[1]_net_1 ), .Y(ADD_26x26_fast_I230_Y_0));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I242_Y (.A(\state[1]_net_1 ), .B(
        LED_FB[5]), .C(N646), .Y(\un1_integ[12] ));
    DFN1E0C0 \integ[11]  (.D(\un1_integ[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(LED_FB[4]));
    DFN1E0C0 \integ[16]  (.D(\un1_integ[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[16]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_1 (.A(
        ADD_26x26_fast_I211_un1_Y_0), .B(N516), .C(
        ADD_26x26_fast_I211_Y_0), .Y(ADD_26x26_fast_I211_Y_1));
    NOR2A \state_RNIV9T8[1]  (.A(\state[1]_net_1 ), .B(avg_old[3]), .Y(
        \un18_next_int_m[3] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I189_Y (.A(N524), .B(N539), .C(
        N523), .Y(N640));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I254_Y_0 (.A(\integ[24]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I254_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I163_Y (.A(I163_un1_Y), .B(N489), 
        .Y(N543));
    AO1 un1_integ_0_0_ADD_26x26_fast_I96_Y (.A(N418), .B(N415), .C(
        N414), .Y(N467));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I207_un1_Y (.A(N524), .B(N508), 
        .C(N539), .Y(I207_un1_Y));
    OR2 \state_RNI7MH81[1]  (.A(\inf_abs0_m[2] ), .B(
        \un18_next_int_m[2] ), .Y(\un1_next_int[2] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I2_G0N (.A(\un1_next_int[2] ), 
        .B(average[2]), .Y(N323));
    OR2 un1_integ_0_0_ADD_26x26_fast_I114_Y (.A(I114_un1_Y), .B(N432), 
        .Y(N485));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I147_Y (.A(N470), .B(N478), .Y(
        N524));
    DFN1E0C0 \integ[9]  (.D(\un1_integ[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(LED_FB[2]));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I235_Y (.A(
        ADD_26x26_fast_I235_Y_0), .B(N541), .Y(\un1_integ[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I212_Y_0 (.A(
        ADD_26x26_fast_I212_un1_Y_0), .B(N518), .C(N517), .Y(
        ADD_26x26_fast_I212_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I63_Y (.A(N336), .B(N333), .Y(
        N431));
    NOR2B \state_1_RNI7BKV[0]  (.A(avg_new[0]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[0] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I118_Y (.A(N440), .B(N437), .C(
        N436), .Y(N489));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I237_Y (.A(\un1_next_int[7] ), 
        .B(LED_FB[0]), .C(N537), .Y(\un1_integ[7] ));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I133_Y (.A(N407), .B(N403), .C(
        N464), .Y(N510));
    OA1B un1_integ_0_0_ADD_26x26_fast_I30_Y (.A(\integ[21]_net_1 ), .B(
        \integ[22]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N398));
    DFN1E0C0 \integ[22]  (.D(\un1_integ[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[22]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I43_Y (.A(\integ[15]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_1[0]_net_1 ), .Y(N411));
    NOR2A \state_RNI5GT8[1]  (.A(\state[1]_net_1 ), .B(avg_old[9]), .Y(
        \un18_next_int_m[9] ));
    DFN1C0 \integ[1]  (.D(ADD_26x26_fast_I231_Y), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\integ[1]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I35_Y (.A(\integ[19]_net_1 ), .B(
        \integ[20]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N403));
    OR2 \state_RNIBQH81[1]  (.A(\un18_next_int_m[4] ), .B(
        \inf_abs0_m[4] ), .Y(\un1_next_int[4] ));
    DFN1C0 \state_0[0]  (.D(\state_RNI3U7Q[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_0[0]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I204_Y_1 (.A(
        ADD_26x26_fast_I204_Y_0), .B(N398), .Y(ADD_26x26_fast_I204_Y_1)
        );
    NOR2B un1_integ_0_0_ADD_26x26_fast_I53_Y (.A(N351), .B(N348), .Y(
        N421));
    AO1 un1_integ_0_0_ADD_26x26_fast_I160_Y (.A(N484), .B(N491), .C(
        N483), .Y(N537));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I91_Y (.A(N413), .B(N409), .Y(
        N462));
    AX1D un1_integ_0_0_ADD_26x26_fast_I250_Y (.A(I178_un1_Y), .B(
        ADD_26x26_fast_I209_Y_1), .C(ADD_26x26_fast_I250_Y_0), .Y(
        \un1_integ[20] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I240_Y_0 (.A(\inf_abs0_m[10] ), 
        .B(\un18_next_int_m[10] ), .C(LED_FB[3]), .Y(
        ADD_26x26_fast_I240_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_0 (.A(N467), .B(N460), .C(
        N459), .Y(ADD_26x26_fast_I210_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I71_Y (.A(average[2]), .B(
        \un1_next_int[2] ), .C(N321), .Y(N439));
    DFN1E0C0 \integ[20]  (.D(\un1_integ[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[20]_net_1 ));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I244_Y (.A(\state_0[0]_net_1 ), 
        .B(LED_FB[7]), .C(N640), .Y(\un1_integ[14] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I207_Y_1 (.A(N404), .B(N400), .C(
        N461), .Y(ADD_26x26_fast_I207_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I106_Y (.A(N428), .B(N425), .C(
        N424), .Y(N477));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_1 (.A(
        ADD_26x26_fast_I208_un1_Y_0), .B(N541), .C(
        ADD_26x26_fast_I208_Y_0), .Y(ADD_26x26_fast_I208_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I102_Y (.A(N424), .B(N421), .C(
        N420), .Y(N473));
    AX1D un1_integ_0_0_ADD_26x26_fast_I251_Y (.A(I176_un1_Y), .B(
        ADD_26x26_fast_I208_Y_1), .C(ADD_26x26_fast_I251_Y_0), .Y(
        \un1_integ[21] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I121_un1_Y (.A(N441), .B(
        \un1_next_int[0] ), .Y(I121_un1_Y));
    DFN1E0C0 \integ[18]  (.D(\un1_integ[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[18]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I4_P0N (.A(average[4]), .B(
        \un1_next_int[4] ), .Y(N330));
    AO1 un1_integ_0_0_ADD_26x26_fast_I144_Y (.A(N475), .B(N468), .C(
        N467), .Y(N521));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I139_Y (.A(N462), .B(N470), .Y(
        N516));
    OR2 \state_RNINB1R[0]  (.A(\inf_abs0_m[11] ), .B(
        \un18_next_int_m[11] ), .Y(\state_RNINB1R[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_0 (.A(N465), .B(N458), .C(
        N457), .Y(ADD_26x26_fast_I209_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I148_Y (.A(N479), .B(N472), .C(
        N471), .Y(N525));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I60_Y (.A(N335), .B(LED_FB[0]), 
        .C(\un1_next_int[7] ), .Y(N428));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y (.A(
        ADD_26x26_fast_I232_Y_0), .B(N493), .Y(ADD_26x26_fast_I232_Y));
    OR3 un1_integ_0_0_ADD_26x26_fast_I204_Y_2 (.A(N406), .B(N402), .C(
        ADD_26x26_fast_I204_Y_1), .Y(ADD_26x26_fast_I204_Y_2));
    DFN1C0 \state[1]  (.D(\state_RNO_3[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[1]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I9_G0N (.A(\un1_next_int[9] ), 
        .B(LED_FB[2]), .Y(N344));
    OA1B un1_integ_0_0_ADD_26x26_fast_I40_Y (.A(\integ[16]_net_1 ), .B(
        \integ[17]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N408));
    OA1 un1_integ_0_0_ADD_26x26_fast_I65_Y (.A(average[4]), .B(
        \un1_next_int[4] ), .C(N333), .Y(N433));
    AO1 un1_integ_0_0_ADD_26x26_fast_I188_Y (.A(N522), .B(N537), .C(
        N521), .Y(N637));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I178_un1_Y (.A(N512), .B(N527), 
        .Y(I178_un1_Y));
    AO1B un1_integ_0_0_ADD_26x26_fast_I45_Y (.A(LED_FB[7]), .B(
        \integ[15]_net_1 ), .C(\state_1[0]_net_1 ), .Y(N413));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I137_Y (.A(N460), .B(N468), .Y(
        N514));
    OR2 un1_integ_0_0_ADD_26x26_fast_I3_P0N (.A(average[3]), .B(
        \un1_next_int[3] ), .Y(N327));
    AO1 un1_integ_0_0_ADD_26x26_fast_I50_Y (.A(N350), .B(N354), .C(
        N353), .Y(N418));
    AO1 un1_integ_0_0_ADD_26x26_fast_I204_Y_3 (.A(N502), .B(N517), .C(
        ADD_26x26_fast_I204_Y_2), .Y(ADD_26x26_fast_I204_Y_3));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I74_un1_Y (.A(N318), .B(
        \un1_next_int[0] ), .Y(I74_un1_Y));
    OA1B un1_integ_0_0_ADD_26x26_fast_I36_Y (.A(\integ[19]_net_1 ), .B(
        \integ[18]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N404));
    OR2 un1_integ_0_0_ADD_26x26_fast_I0_P0N (.A(\integ[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(N318));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I55_Y (.A(N348), .B(N345), .Y(
        N423));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I205_un1_Y (.A(
        ADD_26x26_fast_I205_un1_Y_0), .B(N658), .Y(I205_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I163_un1_Y (.A(N490), .B(
        \un1_next_int[0] ), .Y(I163_un1_Y));
    OR2 \state_RNIJ2I81[1]  (.A(\un18_next_int_m[8] ), .B(
        \inf_abs0_m[8] ), .Y(\un1_next_int[8] ));
    MX2 \un1_integ_0_0_LED_6[4]  (.A(N_54), .B(N_62), .S(choose[1]), 
        .Y(N_70));
    OR3 un1_integ_0_0_ADD_26x26_fast_I206_Y_1 (.A(N398), .B(N402), .C(
        N459), .Y(ADD_26x26_fast_I206_Y_1));
    OA1 un1_integ_0_0_ADD_26x26_fast_I5_G0N (.A(\un18_next_int_m[5] ), 
        .B(\inf_abs0_m[5] ), .C(average[5]), .Y(N332));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I114_un1_Y (.A(N436), .B(N433), 
        .Y(I114_un1_Y));
    DFN1E0C0 \integ[7]  (.D(\un1_integ[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(LED_FB[0]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_2 (.A(N508), .B(N523), .C(
        ADD_26x26_fast_I207_Y_1), .Y(ADD_26x26_fast_I207_Y_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I4_G0N (.A(\un1_next_int[4] ), 
        .B(average[4]), .Y(N329));
    OR2 un1_integ_0_0_ADD_26x26_fast_I195_Y (.A(I195_un1_Y), .B(N535), 
        .Y(N658));
    NOR2B \state_1_RNICGKV[0]  (.A(avg_new[5]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[5] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y (.A(
        ADD_26x26_fast_I234_Y_0), .B(N543), .Y(ADD_26x26_fast_I234_Y));
    OR3 un1_integ_0_0_ADD_26x26_fast_I205_Y_2 (.A(N400), .B(
        ADD_26x26_fast_I205_Y_0), .C(N457), .Y(ADD_26x26_fast_I205_Y_2)
        );
    NOR2B un1_integ_0_0_ADD_26x26_fast_I162_un1_Y (.A(N488), .B(N442), 
        .Y(I162_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I240_Y (.A(N531), .B(I193_un1_Y), 
        .C(ADD_26x26_fast_I240_Y_0), .Y(\un1_integ[10] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I156_Y (.A(N487), .B(N480), .C(
        N479), .Y(N533));
    DFN1E0C0 \integ[8]  (.D(\un1_integ[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(LED_FB[1]));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I251_Y_0 (.A(\integ[21]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I251_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I152_Y (.A(I152_un1_Y), .B(N475), 
        .Y(N529));
    OR2 un1_integ_0_0_ADD_26x26_fast_I9_P0N (.A(\un1_next_int[9] ), .B(
        LED_FB[2]), .Y(N345));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I208_un1_Y_0 (.A(N510), .B(N526)
        , .Y(ADD_26x26_fast_I208_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I191_Y (.A(N528), .B(N543), .C(
        N527), .Y(N646));
    AO1B un1_integ_0_0_ADD_26x26_fast_I31_Y (.A(\integ[21]_net_1 ), .B(
        \integ[22]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N399));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I206_un1_Y (.A(N522), .B(N506), 
        .C(N537), .Y(I206_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I235_Y_0 (.A(
        \un18_next_int_m[5] ), .B(\inf_abs0_m[5] ), .C(average[5]), .Y(
        ADD_26x26_fast_I235_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I241_Y (.A(N529), .B(I192_un1_Y), 
        .C(ADD_26x26_fast_I241_Y_0), .Y(\un1_integ[11] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I11_P0N (.A(
        \state_RNINB1R[0]_net_1 ), .B(LED_FB[4]), .Y(N351));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I243_Y_0 (.A(LED_FB[6]), .B(
        \state[0]_net_1 ), .Y(ADD_26x26_fast_I243_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I105_Y (.A(N423), .B(N427), .Y(
        N476));
    AO1 un1_integ_0_0_ADD_26x26_fast_I213_Y_0 (.A(
        ADD_26x26_fast_I213_un1_Y_0), .B(N520), .C(N519), .Y(
        ADD_26x26_fast_I213_Y_0));
    OR2 \state_RNIFUH81[1]  (.A(\inf_abs0_m[6] ), .B(
        \un18_next_int_m[6] ), .Y(\un1_next_int[6] ));
    NOR2A \state_RNI2DT8[1]  (.A(\state[1]_net_1 ), .B(avg_old[6]), .Y(
        \un18_next_int_m[6] ));
    NOR2B \state_RNI3U7Q[0]  (.A(avg_done), .B(calc_avg), .Y(
        \state_RNI3U7Q[0]_net_1 ));
    NOR2A \state_RNIU8T8[1]  (.A(\state[1]_net_1 ), .B(avg_old[2]), .Y(
        \un18_next_int_m[2] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I101_Y (.A(N419), .B(N423), .Y(
        N472));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I66_Y (.A(N326), .B(average[4]), 
        .C(\un1_next_int[4] ), .Y(N434));
    AX1D un1_integ_0_0_ADD_26x26_fast_I248_Y (.A(I182_un1_Y), .B(
        ADD_26x26_fast_I211_Y_1), .C(ADD_26x26_fast_I248_Y_0), .Y(
        \un1_integ[18] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I99_Y (.A(N417), .B(N421), .Y(
        N470));
    OR2 un1_integ_0_0_ADD_26x26_fast_I92_Y (.A(N414), .B(N410), .Y(
        N463));
    AO1 un1_integ_0_0_ADD_26x26_fast_I72_Y (.A(N317), .B(N321), .C(
        N320), .Y(N440));
    OR2A un1_integ_0_0_ADD_26x26_fast_I13_P0N (.A(\state[0]_net_1 ), 
        .B(LED_FB[6]), .Y(N357));
    NOR2B \state_1_RNIDHKV[0]  (.A(avg_new[6]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[6] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I46_Y (.A(LED_FB[7]), .B(
        LED_FB[6]), .C(\state_1[0]_net_1 ), .Y(N414));
    OR2 \state_RNI5F211[0]  (.A(\inf_abs0_m[9] ), .B(
        \un18_next_int_m[9] ), .Y(\un1_next_int[9] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I116_Y (.A(N438), .B(N435), .C(
        N434), .Y(N487));
    NOR2A \state_RNI3ET8[1]  (.A(\state[1]_net_1 ), .B(avg_old[7]), .Y(
        \un18_next_int_m[7] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I112_Y (.A(I112_un1_Y), .B(N430), 
        .Y(N483));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I8_G0N (.A(\un1_next_int[8] ), 
        .B(LED_FB[1]), .Y(N341));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I213_un1_Y_0 (.A(N482), .B(N490)
        , .C(\un1_next_int[0] ), .Y(ADD_26x26_fast_I213_un1_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y_0 (.A(average[4]), .B(
        \un1_next_int[4] ), .Y(ADD_26x26_fast_I234_Y_0));
    
endmodule


module error_sr_13s_5s_1(
       cur_vd,
       avg_new,
       avg_old,
       avg_enable,
       avg_enable_1,
       avg_enable_0,
       n_rst_c,
       clk_c
    );
input  [11:0] cur_vd;
output [11:0] avg_new;
output [11:0] avg_old;
input  avg_enable;
input  avg_enable_1;
input  avg_enable_0;
input  n_rst_c;
input  clk_c;

    wire \sr_3_[0]_net_1 , \sr_3_[1]_net_1 , \sr_3_[2]_net_1 , 
        \sr_3_[3]_net_1 , \sr_3_[4]_net_1 , \sr_3_[5]_net_1 , 
        \sr_3_[6]_net_1 , \sr_3_[7]_net_1 , \sr_3_[8]_net_1 , 
        \sr_3_[9]_net_1 , \sr_3_[10]_net_1 , \sr_3_[11]_net_1 , 
        \sr_2_[0]_net_1 , \sr_2_[1]_net_1 , \sr_2_[2]_net_1 , 
        \sr_2_[3]_net_1 , \sr_2_[4]_net_1 , \sr_2_[5]_net_1 , 
        \sr_2_[6]_net_1 , \sr_2_[7]_net_1 , \sr_2_[8]_net_1 , 
        \sr_2_[9]_net_1 , \sr_2_[10]_net_1 , \sr_2_[11]_net_1 , 
        \sr_1_[0]_net_1 , \sr_1_[1]_net_1 , \sr_1_[2]_net_1 , 
        \sr_1_[3]_net_1 , \sr_1_[4]_net_1 , \sr_1_[5]_net_1 , 
        \sr_1_[6]_net_1 , \sr_1_[7]_net_1 , \sr_1_[8]_net_1 , 
        \sr_1_[9]_net_1 , \sr_1_[10]_net_1 , \sr_1_[11]_net_1 , GND, 
        VCC;
    
    DFN1E1C0 \sr_1_[11]  (.D(avg_new[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[11]_net_1 ));
    DFN1E1C0 \sr_3_[3]  (.D(\sr_2_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[3]_net_1 ));
    DFN1E1C0 \sr_4_[4]  (.D(\sr_3_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[4]));
    DFN1E1C0 \sr_0_[10]  (.D(cur_vd[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(avg_new[10]));
    DFN1E1C0 \sr_4_[8]  (.D(\sr_3_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[8]));
    DFN1E1C0 \sr_4_[0]  (.D(\sr_3_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[0]));
    DFN1E1C0 \sr_1_[2]  (.D(avg_new[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[2]_net_1 ));
    DFN1E1C0 \sr_0_[2]  (.D(cur_vd[2]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[2]));
    DFN1E1C0 \sr_2_[2]  (.D(\sr_1_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[2]_net_1 ));
    DFN1E1C0 \sr_0_[11]  (.D(cur_vd[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(avg_new[11]));
    DFN1E1C0 \sr_1_[3]  (.D(avg_new[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[3]_net_1 ));
    DFN1E1C0 \sr_0_[3]  (.D(cur_vd[3]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[3]));
    DFN1E1C0 \sr_1_[10]  (.D(avg_new[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[10]_net_1 ));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \sr_4_[10]  (.D(\sr_3_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[10]));
    DFN1E1C0 \sr_3_[11]  (.D(\sr_2_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[11]_net_1 ));
    DFN1E1C0 \sr_2_[3]  (.D(\sr_1_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[3]_net_1 ));
    DFN1E1C0 \sr_3_[6]  (.D(\sr_2_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(\sr_3_[6]_net_1 ));
    DFN1E1C0 \sr_3_[1]  (.D(\sr_2_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[1]_net_1 ));
    DFN1E1C0 \sr_4_[2]  (.D(\sr_3_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[2]));
    DFN1E1C0 \sr_1_[6]  (.D(avg_new[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[6]_net_1 ));
    DFN1E1C0 \sr_4_[3]  (.D(\sr_3_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[3]));
    DFN1E1C0 \sr_0_[6]  (.D(cur_vd[6]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[6]));
    DFN1E1C0 \sr_3_[9]  (.D(\sr_2_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(\sr_3_[9]_net_1 ));
    DFN1E1C0 \sr_1_[1]  (.D(avg_new[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[1]_net_1 ));
    DFN1E1C0 \sr_0_[1]  (.D(cur_vd[1]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[1]));
    DFN1E1C0 \sr_2_[6]  (.D(\sr_1_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[6]_net_1 ));
    DFN1E1C0 \sr_2_[1]  (.D(\sr_1_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[1]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1C0 \sr_3_[5]  (.D(\sr_2_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(\sr_3_[5]_net_1 ));
    DFN1E1C0 \sr_3_[7]  (.D(\sr_2_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(\sr_3_[7]_net_1 ));
    DFN1E1C0 \sr_1_[9]  (.D(avg_new[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(\sr_1_[9]_net_1 ));
    DFN1E1C0 \sr_0_[9]  (.D(cur_vd[9]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[9]));
    DFN1E1C0 \sr_2_[11]  (.D(\sr_1_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(\sr_2_[11]_net_1 ));
    DFN1E1C0 \sr_4_[6]  (.D(\sr_3_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[6]));
    DFN1E1C0 \sr_2_[9]  (.D(\sr_1_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[9]_net_1 ));
    DFN1E1C0 \sr_4_[11]  (.D(\sr_3_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[11]));
    DFN1E1C0 \sr_4_[1]  (.D(\sr_3_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[1]));
    DFN1E1C0 \sr_3_[4]  (.D(\sr_2_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(\sr_3_[4]_net_1 ));
    DFN1E1C0 \sr_1_[5]  (.D(avg_new[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[5]_net_1 ));
    DFN1E1C0 \sr_0_[5]  (.D(cur_vd[5]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[5]));
    DFN1E1C0 \sr_1_[7]  (.D(avg_new[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(\sr_1_[7]_net_1 ));
    DFN1E1C0 \sr_0_[7]  (.D(cur_vd[7]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[7]));
    DFN1E1C0 \sr_3_[8]  (.D(\sr_2_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(\sr_3_[8]_net_1 ));
    DFN1E1C0 \sr_3_[0]  (.D(\sr_2_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[0]_net_1 ));
    DFN1E1C0 \sr_2_[5]  (.D(\sr_1_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[5]_net_1 ));
    DFN1E1C0 \sr_2_[7]  (.D(\sr_1_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[7]_net_1 ));
    DFN1E1C0 \sr_4_[9]  (.D(\sr_3_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[9]));
    DFN1E1C0 \sr_1_[4]  (.D(avg_new[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[4]_net_1 ));
    DFN1E1C0 \sr_0_[4]  (.D(cur_vd[4]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[4]));
    DFN1E1C0 \sr_1_[8]  (.D(avg_new[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(\sr_1_[8]_net_1 ));
    DFN1E1C0 \sr_1_[0]  (.D(avg_new[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[0]_net_1 ));
    DFN1E1C0 \sr_2_[4]  (.D(\sr_1_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[4]_net_1 ));
    DFN1E1C0 \sr_0_[8]  (.D(cur_vd[8]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[8]));
    DFN1E1C0 \sr_0_[0]  (.D(cur_vd[0]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[0]));
    DFN1E1C0 \sr_4_[5]  (.D(\sr_3_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[5]));
    DFN1E1C0 \sr_2_[8]  (.D(\sr_1_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[8]_net_1 ));
    DFN1E1C0 \sr_2_[0]  (.D(\sr_1_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[0]_net_1 ));
    DFN1E1C0 \sr_4_[7]  (.D(\sr_3_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[7]));
    DFN1E1C0 \sr_3_[10]  (.D(\sr_2_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[10]_net_1 ));
    DFN1E1C0 \sr_3_[2]  (.D(\sr_2_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[2]_net_1 ));
    DFN1E1C0 \sr_2_[10]  (.D(\sr_1_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(\sr_2_[10]_net_1 ));
    
endmodule


module error_sr_13s_64s_1(
       sr_old,
       sr_new,
       cur_error,
       sr_prev,
       sr_old_0_0,
       sr_new_0_0,
       sr_new_1_0,
       int_enable_11,
       int_enable_29,
       int_enable_19,
       int_enable_8,
       int_enable_4,
       int_enable_28,
       int_enable_17,
       int_enable_26,
       int_enable_9,
       int_enable_18,
       int_enable_21,
       int_enable_20,
       int_enable_27,
       int_enable_31,
       int_enable_30,
       int_enable_5,
       int_enable_3,
       int_enable_2,
       int_enable_14,
       int_enable_13,
       int_enable_23,
       int_enable_12,
       int_enable_32,
       int_enable_1,
       int_enable_7,
       int_enable_6,
       int_enable_22,
       int_enable_16,
       int_enable_15,
       int_enable_10,
       int_enable_25,
       int_enable_24,
       int_enable_33,
       int_enable,
       int_enable_0,
       n_rst_c,
       clk_c
    );
output [12:0] sr_old;
output [12:0] sr_new;
input  [12:0] cur_error;
output [12:0] sr_prev;
output sr_old_0_0;
output sr_new_0_0;
output sr_new_1_0;
input  int_enable_11;
input  int_enable_29;
input  int_enable_19;
input  int_enable_8;
input  int_enable_4;
input  int_enable_28;
input  int_enable_17;
input  int_enable_26;
input  int_enable_9;
input  int_enable_18;
input  int_enable_21;
input  int_enable_20;
input  int_enable_27;
input  int_enable_31;
input  int_enable_30;
input  int_enable_5;
input  int_enable_3;
input  int_enable_2;
input  int_enable_14;
input  int_enable_13;
input  int_enable_23;
input  int_enable_12;
input  int_enable_32;
input  int_enable_1;
input  int_enable_7;
input  int_enable_6;
input  int_enable_22;
input  int_enable_16;
input  int_enable_15;
input  int_enable_10;
input  int_enable_25;
input  int_enable_24;
input  int_enable_33;
input  int_enable;
input  int_enable_0;
input  n_rst_c;
input  clk_c;

    wire \sr_62_[12]_net_1 , \sr_9_[0]_net_1 , \sr_8_[0]_net_1 , 
        \sr_9_[1]_net_1 , \sr_8_[1]_net_1 , \sr_9_[2]_net_1 , 
        \sr_8_[2]_net_1 , \sr_9_[3]_net_1 , \sr_8_[3]_net_1 , 
        \sr_9_[4]_net_1 , \sr_8_[4]_net_1 , \sr_9_[5]_net_1 , 
        \sr_8_[5]_net_1 , \sr_9_[6]_net_1 , \sr_8_[6]_net_1 , 
        \sr_9_[7]_net_1 , \sr_8_[7]_net_1 , \sr_9_[8]_net_1 , 
        \sr_8_[8]_net_1 , \sr_9_[9]_net_1 , \sr_8_[9]_net_1 , 
        \sr_9_[10]_net_1 , \sr_8_[10]_net_1 , \sr_9_[11]_net_1 , 
        \sr_8_[11]_net_1 , \sr_9_[12]_net_1 , \sr_8_[12]_net_1 , 
        \sr_7_[0]_net_1 , \sr_7_[1]_net_1 , \sr_7_[2]_net_1 , 
        \sr_7_[3]_net_1 , \sr_7_[4]_net_1 , \sr_7_[5]_net_1 , 
        \sr_7_[6]_net_1 , \sr_7_[7]_net_1 , \sr_7_[8]_net_1 , 
        \sr_7_[9]_net_1 , \sr_7_[10]_net_1 , \sr_7_[11]_net_1 , 
        \sr_7_[12]_net_1 , \sr_6_[0]_net_1 , \sr_6_[1]_net_1 , 
        \sr_6_[2]_net_1 , \sr_6_[3]_net_1 , \sr_6_[4]_net_1 , 
        \sr_6_[5]_net_1 , \sr_6_[6]_net_1 , \sr_6_[7]_net_1 , 
        \sr_6_[8]_net_1 , \sr_6_[9]_net_1 , \sr_6_[10]_net_1 , 
        \sr_6_[11]_net_1 , \sr_6_[12]_net_1 , \sr_5_[0]_net_1 , 
        \sr_5_[1]_net_1 , \sr_5_[2]_net_1 , \sr_5_[3]_net_1 , 
        \sr_5_[4]_net_1 , \sr_5_[5]_net_1 , \sr_5_[6]_net_1 , 
        \sr_5_[7]_net_1 , \sr_5_[8]_net_1 , \sr_5_[9]_net_1 , 
        \sr_5_[10]_net_1 , \sr_5_[11]_net_1 , \sr_5_[12]_net_1 , 
        \sr_4_[0]_net_1 , \sr_4_[1]_net_1 , \sr_4_[2]_net_1 , 
        \sr_4_[3]_net_1 , \sr_4_[4]_net_1 , \sr_4_[5]_net_1 , 
        \sr_4_[6]_net_1 , \sr_4_[7]_net_1 , \sr_4_[8]_net_1 , 
        \sr_4_[9]_net_1 , \sr_4_[10]_net_1 , \sr_4_[11]_net_1 , 
        \sr_4_[12]_net_1 , \sr_3_[0]_net_1 , \sr_3_[1]_net_1 , 
        \sr_3_[2]_net_1 , \sr_3_[3]_net_1 , \sr_3_[4]_net_1 , 
        \sr_3_[5]_net_1 , \sr_3_[6]_net_1 , \sr_3_[7]_net_1 , 
        \sr_3_[8]_net_1 , \sr_3_[9]_net_1 , \sr_3_[10]_net_1 , 
        \sr_3_[11]_net_1 , \sr_3_[12]_net_1 , \sr_2_[0]_net_1 , 
        \sr_2_[1]_net_1 , \sr_2_[2]_net_1 , \sr_2_[3]_net_1 , 
        \sr_2_[4]_net_1 , \sr_2_[5]_net_1 , \sr_2_[6]_net_1 , 
        \sr_2_[7]_net_1 , \sr_2_[8]_net_1 , \sr_2_[9]_net_1 , 
        \sr_2_[10]_net_1 , \sr_2_[11]_net_1 , \sr_2_[12]_net_1 , 
        \sr_24_[0]_net_1 , \sr_23_[0]_net_1 , \sr_24_[1]_net_1 , 
        \sr_23_[1]_net_1 , \sr_24_[2]_net_1 , \sr_23_[2]_net_1 , 
        \sr_24_[3]_net_1 , \sr_23_[3]_net_1 , \sr_24_[4]_net_1 , 
        \sr_23_[4]_net_1 , \sr_24_[5]_net_1 , \sr_23_[5]_net_1 , 
        \sr_24_[6]_net_1 , \sr_23_[6]_net_1 , \sr_24_[7]_net_1 , 
        \sr_23_[7]_net_1 , \sr_24_[8]_net_1 , \sr_23_[8]_net_1 , 
        \sr_24_[9]_net_1 , \sr_23_[9]_net_1 , \sr_24_[10]_net_1 , 
        \sr_23_[10]_net_1 , \sr_24_[11]_net_1 , \sr_23_[11]_net_1 , 
        \sr_24_[12]_net_1 , \sr_23_[12]_net_1 , \sr_22_[0]_net_1 , 
        \sr_22_[1]_net_1 , \sr_22_[2]_net_1 , \sr_22_[3]_net_1 , 
        \sr_22_[4]_net_1 , \sr_22_[5]_net_1 , \sr_22_[6]_net_1 , 
        \sr_22_[7]_net_1 , \sr_22_[8]_net_1 , \sr_22_[9]_net_1 , 
        \sr_22_[10]_net_1 , \sr_22_[11]_net_1 , \sr_22_[12]_net_1 , 
        \sr_21_[0]_net_1 , \sr_21_[1]_net_1 , \sr_21_[2]_net_1 , 
        \sr_21_[3]_net_1 , \sr_21_[4]_net_1 , \sr_21_[5]_net_1 , 
        \sr_21_[6]_net_1 , \sr_21_[7]_net_1 , \sr_21_[8]_net_1 , 
        \sr_21_[9]_net_1 , \sr_21_[10]_net_1 , \sr_21_[11]_net_1 , 
        \sr_21_[12]_net_1 , \sr_20_[0]_net_1 , \sr_20_[1]_net_1 , 
        \sr_20_[2]_net_1 , \sr_20_[3]_net_1 , \sr_20_[4]_net_1 , 
        \sr_20_[5]_net_1 , \sr_20_[6]_net_1 , \sr_20_[7]_net_1 , 
        \sr_20_[8]_net_1 , \sr_20_[9]_net_1 , \sr_20_[10]_net_1 , 
        \sr_20_[11]_net_1 , \sr_20_[12]_net_1 , \sr_19_[0]_net_1 , 
        \sr_19_[1]_net_1 , \sr_19_[2]_net_1 , \sr_19_[3]_net_1 , 
        \sr_19_[4]_net_1 , \sr_19_[5]_net_1 , \sr_19_[6]_net_1 , 
        \sr_19_[7]_net_1 , \sr_19_[8]_net_1 , \sr_19_[9]_net_1 , 
        \sr_19_[10]_net_1 , \sr_19_[11]_net_1 , \sr_19_[12]_net_1 , 
        \sr_18_[0]_net_1 , \sr_18_[1]_net_1 , \sr_18_[2]_net_1 , 
        \sr_18_[3]_net_1 , \sr_18_[4]_net_1 , \sr_18_[5]_net_1 , 
        \sr_18_[6]_net_1 , \sr_18_[7]_net_1 , \sr_18_[8]_net_1 , 
        \sr_18_[9]_net_1 , \sr_18_[10]_net_1 , \sr_18_[11]_net_1 , 
        \sr_18_[12]_net_1 , \sr_17_[0]_net_1 , \sr_17_[1]_net_1 , 
        \sr_17_[2]_net_1 , \sr_17_[3]_net_1 , \sr_17_[4]_net_1 , 
        \sr_17_[5]_net_1 , \sr_17_[6]_net_1 , \sr_17_[7]_net_1 , 
        \sr_17_[8]_net_1 , \sr_17_[9]_net_1 , \sr_17_[10]_net_1 , 
        \sr_17_[11]_net_1 , \sr_17_[12]_net_1 , \sr_16_[0]_net_1 , 
        \sr_16_[1]_net_1 , \sr_16_[2]_net_1 , \sr_16_[3]_net_1 , 
        \sr_16_[4]_net_1 , \sr_16_[5]_net_1 , \sr_16_[6]_net_1 , 
        \sr_16_[7]_net_1 , \sr_16_[8]_net_1 , \sr_16_[9]_net_1 , 
        \sr_16_[10]_net_1 , \sr_16_[11]_net_1 , \sr_16_[12]_net_1 , 
        \sr_15_[0]_net_1 , \sr_15_[1]_net_1 , \sr_15_[2]_net_1 , 
        \sr_15_[3]_net_1 , \sr_15_[4]_net_1 , \sr_15_[5]_net_1 , 
        \sr_15_[6]_net_1 , \sr_15_[7]_net_1 , \sr_15_[8]_net_1 , 
        \sr_15_[9]_net_1 , \sr_15_[10]_net_1 , \sr_15_[11]_net_1 , 
        \sr_15_[12]_net_1 , \sr_14_[0]_net_1 , \sr_14_[1]_net_1 , 
        \sr_14_[2]_net_1 , \sr_14_[3]_net_1 , \sr_14_[4]_net_1 , 
        \sr_14_[5]_net_1 , \sr_14_[6]_net_1 , \sr_14_[7]_net_1 , 
        \sr_14_[8]_net_1 , \sr_14_[9]_net_1 , \sr_14_[10]_net_1 , 
        \sr_14_[11]_net_1 , \sr_14_[12]_net_1 , \sr_13_[0]_net_1 , 
        \sr_13_[1]_net_1 , \sr_13_[2]_net_1 , \sr_13_[3]_net_1 , 
        \sr_13_[4]_net_1 , \sr_13_[5]_net_1 , \sr_13_[6]_net_1 , 
        \sr_13_[7]_net_1 , \sr_13_[8]_net_1 , \sr_13_[9]_net_1 , 
        \sr_13_[10]_net_1 , \sr_13_[11]_net_1 , \sr_13_[12]_net_1 , 
        \sr_12_[0]_net_1 , \sr_12_[1]_net_1 , \sr_12_[2]_net_1 , 
        \sr_12_[3]_net_1 , \sr_12_[4]_net_1 , \sr_12_[5]_net_1 , 
        \sr_12_[6]_net_1 , \sr_12_[7]_net_1 , \sr_12_[8]_net_1 , 
        \sr_12_[9]_net_1 , \sr_12_[10]_net_1 , \sr_12_[11]_net_1 , 
        \sr_12_[12]_net_1 , \sr_11_[0]_net_1 , \sr_11_[1]_net_1 , 
        \sr_11_[2]_net_1 , \sr_11_[3]_net_1 , \sr_11_[4]_net_1 , 
        \sr_11_[5]_net_1 , \sr_11_[6]_net_1 , \sr_11_[7]_net_1 , 
        \sr_11_[8]_net_1 , \sr_11_[9]_net_1 , \sr_11_[10]_net_1 , 
        \sr_11_[11]_net_1 , \sr_11_[12]_net_1 , \sr_10_[0]_net_1 , 
        \sr_10_[1]_net_1 , \sr_10_[2]_net_1 , \sr_10_[3]_net_1 , 
        \sr_10_[4]_net_1 , \sr_10_[5]_net_1 , \sr_10_[6]_net_1 , 
        \sr_10_[7]_net_1 , \sr_10_[8]_net_1 , \sr_10_[9]_net_1 , 
        \sr_10_[10]_net_1 , \sr_10_[11]_net_1 , \sr_10_[12]_net_1 , 
        \sr_39_[0]_net_1 , \sr_38_[0]_net_1 , \sr_39_[1]_net_1 , 
        \sr_38_[1]_net_1 , \sr_39_[2]_net_1 , \sr_38_[2]_net_1 , 
        \sr_39_[3]_net_1 , \sr_38_[3]_net_1 , \sr_39_[4]_net_1 , 
        \sr_38_[4]_net_1 , \sr_39_[5]_net_1 , \sr_38_[5]_net_1 , 
        \sr_39_[6]_net_1 , \sr_38_[6]_net_1 , \sr_39_[7]_net_1 , 
        \sr_38_[7]_net_1 , \sr_39_[8]_net_1 , \sr_38_[8]_net_1 , 
        \sr_39_[9]_net_1 , \sr_38_[9]_net_1 , \sr_39_[10]_net_1 , 
        \sr_38_[10]_net_1 , \sr_39_[11]_net_1 , \sr_38_[11]_net_1 , 
        \sr_39_[12]_net_1 , \sr_38_[12]_net_1 , \sr_37_[0]_net_1 , 
        \sr_37_[1]_net_1 , \sr_37_[2]_net_1 , \sr_37_[3]_net_1 , 
        \sr_37_[4]_net_1 , \sr_37_[5]_net_1 , \sr_37_[6]_net_1 , 
        \sr_37_[7]_net_1 , \sr_37_[8]_net_1 , \sr_37_[9]_net_1 , 
        \sr_37_[10]_net_1 , \sr_37_[11]_net_1 , \sr_37_[12]_net_1 , 
        \sr_36_[0]_net_1 , \sr_36_[1]_net_1 , \sr_36_[2]_net_1 , 
        \sr_36_[3]_net_1 , \sr_36_[4]_net_1 , \sr_36_[5]_net_1 , 
        \sr_36_[6]_net_1 , \sr_36_[7]_net_1 , \sr_36_[8]_net_1 , 
        \sr_36_[9]_net_1 , \sr_36_[10]_net_1 , \sr_36_[11]_net_1 , 
        \sr_36_[12]_net_1 , \sr_35_[0]_net_1 , \sr_35_[1]_net_1 , 
        \sr_35_[2]_net_1 , \sr_35_[3]_net_1 , \sr_35_[4]_net_1 , 
        \sr_35_[5]_net_1 , \sr_35_[6]_net_1 , \sr_35_[7]_net_1 , 
        \sr_35_[8]_net_1 , \sr_35_[9]_net_1 , \sr_35_[10]_net_1 , 
        \sr_35_[11]_net_1 , \sr_35_[12]_net_1 , \sr_34_[0]_net_1 , 
        \sr_34_[1]_net_1 , \sr_34_[2]_net_1 , \sr_34_[3]_net_1 , 
        \sr_34_[4]_net_1 , \sr_34_[5]_net_1 , \sr_34_[6]_net_1 , 
        \sr_34_[7]_net_1 , \sr_34_[8]_net_1 , \sr_34_[9]_net_1 , 
        \sr_34_[10]_net_1 , \sr_34_[11]_net_1 , \sr_34_[12]_net_1 , 
        \sr_33_[0]_net_1 , \sr_33_[1]_net_1 , \sr_33_[2]_net_1 , 
        \sr_33_[3]_net_1 , \sr_33_[4]_net_1 , \sr_33_[5]_net_1 , 
        \sr_33_[6]_net_1 , \sr_33_[7]_net_1 , \sr_33_[8]_net_1 , 
        \sr_33_[9]_net_1 , \sr_33_[10]_net_1 , \sr_33_[11]_net_1 , 
        \sr_33_[12]_net_1 , \sr_32_[0]_net_1 , \sr_32_[1]_net_1 , 
        \sr_32_[2]_net_1 , \sr_32_[3]_net_1 , \sr_32_[4]_net_1 , 
        \sr_32_[5]_net_1 , \sr_32_[6]_net_1 , \sr_32_[7]_net_1 , 
        \sr_32_[8]_net_1 , \sr_32_[9]_net_1 , \sr_32_[10]_net_1 , 
        \sr_32_[11]_net_1 , \sr_32_[12]_net_1 , \sr_31_[0]_net_1 , 
        \sr_31_[1]_net_1 , \sr_31_[2]_net_1 , \sr_31_[3]_net_1 , 
        \sr_31_[4]_net_1 , \sr_31_[5]_net_1 , \sr_31_[6]_net_1 , 
        \sr_31_[7]_net_1 , \sr_31_[8]_net_1 , \sr_31_[9]_net_1 , 
        \sr_31_[10]_net_1 , \sr_31_[11]_net_1 , \sr_31_[12]_net_1 , 
        \sr_30_[0]_net_1 , \sr_30_[1]_net_1 , \sr_30_[2]_net_1 , 
        \sr_30_[3]_net_1 , \sr_30_[4]_net_1 , \sr_30_[5]_net_1 , 
        \sr_30_[6]_net_1 , \sr_30_[7]_net_1 , \sr_30_[8]_net_1 , 
        \sr_30_[9]_net_1 , \sr_30_[10]_net_1 , \sr_30_[11]_net_1 , 
        \sr_30_[12]_net_1 , \sr_29_[0]_net_1 , \sr_29_[1]_net_1 , 
        \sr_29_[2]_net_1 , \sr_29_[3]_net_1 , \sr_29_[4]_net_1 , 
        \sr_29_[5]_net_1 , \sr_29_[6]_net_1 , \sr_29_[7]_net_1 , 
        \sr_29_[8]_net_1 , \sr_29_[9]_net_1 , \sr_29_[10]_net_1 , 
        \sr_29_[11]_net_1 , \sr_29_[12]_net_1 , \sr_28_[0]_net_1 , 
        \sr_28_[1]_net_1 , \sr_28_[2]_net_1 , \sr_28_[3]_net_1 , 
        \sr_28_[4]_net_1 , \sr_28_[5]_net_1 , \sr_28_[6]_net_1 , 
        \sr_28_[7]_net_1 , \sr_28_[8]_net_1 , \sr_28_[9]_net_1 , 
        \sr_28_[10]_net_1 , \sr_28_[11]_net_1 , \sr_28_[12]_net_1 , 
        \sr_27_[0]_net_1 , \sr_27_[1]_net_1 , \sr_27_[2]_net_1 , 
        \sr_27_[3]_net_1 , \sr_27_[4]_net_1 , \sr_27_[5]_net_1 , 
        \sr_27_[6]_net_1 , \sr_27_[7]_net_1 , \sr_27_[8]_net_1 , 
        \sr_27_[9]_net_1 , \sr_27_[10]_net_1 , \sr_27_[11]_net_1 , 
        \sr_27_[12]_net_1 , \sr_26_[0]_net_1 , \sr_26_[1]_net_1 , 
        \sr_26_[2]_net_1 , \sr_26_[3]_net_1 , \sr_26_[4]_net_1 , 
        \sr_26_[5]_net_1 , \sr_26_[6]_net_1 , \sr_26_[7]_net_1 , 
        \sr_26_[8]_net_1 , \sr_26_[9]_net_1 , \sr_26_[10]_net_1 , 
        \sr_26_[11]_net_1 , \sr_26_[12]_net_1 , \sr_25_[0]_net_1 , 
        \sr_25_[1]_net_1 , \sr_25_[2]_net_1 , \sr_25_[3]_net_1 , 
        \sr_25_[4]_net_1 , \sr_25_[5]_net_1 , \sr_25_[6]_net_1 , 
        \sr_25_[7]_net_1 , \sr_25_[8]_net_1 , \sr_25_[9]_net_1 , 
        \sr_25_[10]_net_1 , \sr_25_[11]_net_1 , \sr_25_[12]_net_1 , 
        \sr_54_[0]_net_1 , \sr_53_[0]_net_1 , \sr_54_[1]_net_1 , 
        \sr_53_[1]_net_1 , \sr_54_[2]_net_1 , \sr_53_[2]_net_1 , 
        \sr_54_[3]_net_1 , \sr_53_[3]_net_1 , \sr_54_[4]_net_1 , 
        \sr_53_[4]_net_1 , \sr_54_[5]_net_1 , \sr_53_[5]_net_1 , 
        \sr_54_[6]_net_1 , \sr_53_[6]_net_1 , \sr_54_[7]_net_1 , 
        \sr_53_[7]_net_1 , \sr_54_[8]_net_1 , \sr_53_[8]_net_1 , 
        \sr_54_[9]_net_1 , \sr_53_[9]_net_1 , \sr_54_[10]_net_1 , 
        \sr_53_[10]_net_1 , \sr_54_[11]_net_1 , \sr_53_[11]_net_1 , 
        \sr_54_[12]_net_1 , \sr_53_[12]_net_1 , \sr_52_[0]_net_1 , 
        \sr_52_[1]_net_1 , \sr_52_[2]_net_1 , \sr_52_[3]_net_1 , 
        \sr_52_[4]_net_1 , \sr_52_[5]_net_1 , \sr_52_[6]_net_1 , 
        \sr_52_[7]_net_1 , \sr_52_[8]_net_1 , \sr_52_[9]_net_1 , 
        \sr_52_[10]_net_1 , \sr_52_[11]_net_1 , \sr_52_[12]_net_1 , 
        \sr_51_[0]_net_1 , \sr_51_[1]_net_1 , \sr_51_[2]_net_1 , 
        \sr_51_[3]_net_1 , \sr_51_[4]_net_1 , \sr_51_[5]_net_1 , 
        \sr_51_[6]_net_1 , \sr_51_[7]_net_1 , \sr_51_[8]_net_1 , 
        \sr_51_[9]_net_1 , \sr_51_[10]_net_1 , \sr_51_[11]_net_1 , 
        \sr_51_[12]_net_1 , \sr_50_[0]_net_1 , \sr_50_[1]_net_1 , 
        \sr_50_[2]_net_1 , \sr_50_[3]_net_1 , \sr_50_[4]_net_1 , 
        \sr_50_[5]_net_1 , \sr_50_[6]_net_1 , \sr_50_[7]_net_1 , 
        \sr_50_[8]_net_1 , \sr_50_[9]_net_1 , \sr_50_[10]_net_1 , 
        \sr_50_[11]_net_1 , \sr_50_[12]_net_1 , \sr_49_[0]_net_1 , 
        \sr_49_[1]_net_1 , \sr_49_[2]_net_1 , \sr_49_[3]_net_1 , 
        \sr_49_[4]_net_1 , \sr_49_[5]_net_1 , \sr_49_[6]_net_1 , 
        \sr_49_[7]_net_1 , \sr_49_[8]_net_1 , \sr_49_[9]_net_1 , 
        \sr_49_[10]_net_1 , \sr_49_[11]_net_1 , \sr_49_[12]_net_1 , 
        \sr_48_[0]_net_1 , \sr_48_[1]_net_1 , \sr_48_[2]_net_1 , 
        \sr_48_[3]_net_1 , \sr_48_[4]_net_1 , \sr_48_[5]_net_1 , 
        \sr_48_[6]_net_1 , \sr_48_[7]_net_1 , \sr_48_[8]_net_1 , 
        \sr_48_[9]_net_1 , \sr_48_[10]_net_1 , \sr_48_[11]_net_1 , 
        \sr_48_[12]_net_1 , \sr_47_[0]_net_1 , \sr_47_[1]_net_1 , 
        \sr_47_[2]_net_1 , \sr_47_[3]_net_1 , \sr_47_[4]_net_1 , 
        \sr_47_[5]_net_1 , \sr_47_[6]_net_1 , \sr_47_[7]_net_1 , 
        \sr_47_[8]_net_1 , \sr_47_[9]_net_1 , \sr_47_[10]_net_1 , 
        \sr_47_[11]_net_1 , \sr_47_[12]_net_1 , \sr_46_[0]_net_1 , 
        \sr_46_[1]_net_1 , \sr_46_[2]_net_1 , \sr_46_[3]_net_1 , 
        \sr_46_[4]_net_1 , \sr_46_[5]_net_1 , \sr_46_[6]_net_1 , 
        \sr_46_[7]_net_1 , \sr_46_[8]_net_1 , \sr_46_[9]_net_1 , 
        \sr_46_[10]_net_1 , \sr_46_[11]_net_1 , \sr_46_[12]_net_1 , 
        \sr_45_[0]_net_1 , \sr_45_[1]_net_1 , \sr_45_[2]_net_1 , 
        \sr_45_[3]_net_1 , \sr_45_[4]_net_1 , \sr_45_[5]_net_1 , 
        \sr_45_[6]_net_1 , \sr_45_[7]_net_1 , \sr_45_[8]_net_1 , 
        \sr_45_[9]_net_1 , \sr_45_[10]_net_1 , \sr_45_[11]_net_1 , 
        \sr_45_[12]_net_1 , \sr_44_[0]_net_1 , \sr_44_[1]_net_1 , 
        \sr_44_[2]_net_1 , \sr_44_[3]_net_1 , \sr_44_[4]_net_1 , 
        \sr_44_[5]_net_1 , \sr_44_[6]_net_1 , \sr_44_[7]_net_1 , 
        \sr_44_[8]_net_1 , \sr_44_[9]_net_1 , \sr_44_[10]_net_1 , 
        \sr_44_[11]_net_1 , \sr_44_[12]_net_1 , \sr_43_[0]_net_1 , 
        \sr_43_[1]_net_1 , \sr_43_[2]_net_1 , \sr_43_[3]_net_1 , 
        \sr_43_[4]_net_1 , \sr_43_[5]_net_1 , \sr_43_[6]_net_1 , 
        \sr_43_[7]_net_1 , \sr_43_[8]_net_1 , \sr_43_[9]_net_1 , 
        \sr_43_[10]_net_1 , \sr_43_[11]_net_1 , \sr_43_[12]_net_1 , 
        \sr_42_[0]_net_1 , \sr_42_[1]_net_1 , \sr_42_[2]_net_1 , 
        \sr_42_[3]_net_1 , \sr_42_[4]_net_1 , \sr_42_[5]_net_1 , 
        \sr_42_[6]_net_1 , \sr_42_[7]_net_1 , \sr_42_[8]_net_1 , 
        \sr_42_[9]_net_1 , \sr_42_[10]_net_1 , \sr_42_[11]_net_1 , 
        \sr_42_[12]_net_1 , \sr_41_[0]_net_1 , \sr_41_[1]_net_1 , 
        \sr_41_[2]_net_1 , \sr_41_[3]_net_1 , \sr_41_[4]_net_1 , 
        \sr_41_[5]_net_1 , \sr_41_[6]_net_1 , \sr_41_[7]_net_1 , 
        \sr_41_[8]_net_1 , \sr_41_[9]_net_1 , \sr_41_[10]_net_1 , 
        \sr_41_[11]_net_1 , \sr_41_[12]_net_1 , \sr_40_[0]_net_1 , 
        \sr_40_[1]_net_1 , \sr_40_[2]_net_1 , \sr_40_[3]_net_1 , 
        \sr_40_[4]_net_1 , \sr_40_[5]_net_1 , \sr_40_[6]_net_1 , 
        \sr_40_[7]_net_1 , \sr_40_[8]_net_1 , \sr_40_[9]_net_1 , 
        \sr_40_[10]_net_1 , \sr_40_[11]_net_1 , \sr_40_[12]_net_1 , 
        \sr_62_[0]_net_1 , \sr_62_[1]_net_1 , \sr_62_[2]_net_1 , 
        \sr_62_[3]_net_1 , \sr_62_[4]_net_1 , \sr_62_[5]_net_1 , 
        \sr_62_[6]_net_1 , \sr_62_[7]_net_1 , \sr_62_[8]_net_1 , 
        \sr_62_[9]_net_1 , \sr_62_[10]_net_1 , \sr_62_[11]_net_1 , 
        \sr_61_[0]_net_1 , \sr_61_[1]_net_1 , \sr_61_[2]_net_1 , 
        \sr_61_[3]_net_1 , \sr_61_[4]_net_1 , \sr_61_[5]_net_1 , 
        \sr_61_[6]_net_1 , \sr_61_[7]_net_1 , \sr_61_[8]_net_1 , 
        \sr_61_[9]_net_1 , \sr_61_[10]_net_1 , \sr_61_[11]_net_1 , 
        \sr_61_[12]_net_1 , \sr_60_[0]_net_1 , \sr_60_[1]_net_1 , 
        \sr_60_[2]_net_1 , \sr_60_[3]_net_1 , \sr_60_[4]_net_1 , 
        \sr_60_[5]_net_1 , \sr_60_[6]_net_1 , \sr_60_[7]_net_1 , 
        \sr_60_[8]_net_1 , \sr_60_[9]_net_1 , \sr_60_[10]_net_1 , 
        \sr_60_[11]_net_1 , \sr_60_[12]_net_1 , \sr_59_[0]_net_1 , 
        \sr_59_[1]_net_1 , \sr_59_[2]_net_1 , \sr_59_[3]_net_1 , 
        \sr_59_[4]_net_1 , \sr_59_[5]_net_1 , \sr_59_[6]_net_1 , 
        \sr_59_[7]_net_1 , \sr_59_[8]_net_1 , \sr_59_[9]_net_1 , 
        \sr_59_[10]_net_1 , \sr_59_[11]_net_1 , \sr_59_[12]_net_1 , 
        \sr_58_[0]_net_1 , \sr_58_[1]_net_1 , \sr_58_[2]_net_1 , 
        \sr_58_[3]_net_1 , \sr_58_[4]_net_1 , \sr_58_[5]_net_1 , 
        \sr_58_[6]_net_1 , \sr_58_[7]_net_1 , \sr_58_[8]_net_1 , 
        \sr_58_[9]_net_1 , \sr_58_[10]_net_1 , \sr_58_[11]_net_1 , 
        \sr_58_[12]_net_1 , \sr_57_[0]_net_1 , \sr_57_[1]_net_1 , 
        \sr_57_[2]_net_1 , \sr_57_[3]_net_1 , \sr_57_[4]_net_1 , 
        \sr_57_[5]_net_1 , \sr_57_[6]_net_1 , \sr_57_[7]_net_1 , 
        \sr_57_[8]_net_1 , \sr_57_[9]_net_1 , \sr_57_[10]_net_1 , 
        \sr_57_[11]_net_1 , \sr_57_[12]_net_1 , \sr_56_[0]_net_1 , 
        \sr_56_[1]_net_1 , \sr_56_[2]_net_1 , \sr_56_[3]_net_1 , 
        \sr_56_[4]_net_1 , \sr_56_[5]_net_1 , \sr_56_[6]_net_1 , 
        \sr_56_[7]_net_1 , \sr_56_[8]_net_1 , \sr_56_[9]_net_1 , 
        \sr_56_[10]_net_1 , \sr_56_[11]_net_1 , \sr_56_[12]_net_1 , 
        \sr_55_[0]_net_1 , \sr_55_[1]_net_1 , \sr_55_[2]_net_1 , 
        \sr_55_[3]_net_1 , \sr_55_[4]_net_1 , \sr_55_[5]_net_1 , 
        \sr_55_[6]_net_1 , \sr_55_[7]_net_1 , \sr_55_[8]_net_1 , 
        \sr_55_[9]_net_1 , \sr_55_[10]_net_1 , \sr_55_[11]_net_1 , 
        \sr_55_[12]_net_1 , GND, VCC;
    
    DFN1E1C0 \sr_41_[5]  (.D(\sr_40_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_41_[5]_net_1 ));
    DFN1E1C0 \sr_15_[3]  (.D(\sr_14_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_5), .Q(\sr_15_[3]_net_1 ));
    DFN1E1C0 \sr_36_[5]  (.D(\sr_35_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_36_[5]_net_1 ));
    DFN1E1C0 \sr_57_[5]  (.D(\sr_56_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_57_[5]_net_1 ));
    DFN1E1C0 \sr_45_[11]  (.D(\sr_44_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_45_[11]_net_1 ));
    DFN1E1C0 \sr_39_[6]  (.D(\sr_38_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_39_[6]_net_1 ));
    DFN1E1C0 \sr_36_[4]  (.D(\sr_35_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_36_[4]_net_1 ));
    DFN1E1C0 \sr_42_[4]  (.D(\sr_41_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_42_[4]_net_1 ));
    DFN1E1C0 \sr_9_[3]  (.D(\sr_8_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[3]_net_1 ));
    DFN1E1C0 \sr_6_[4]  (.D(\sr_5_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_6_[4]_net_1 ));
    DFN1E1C0 \sr_32_[3]  (.D(\sr_31_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_32_[3]_net_1 ));
    DFN1E1C0 \sr_52_[6]  (.D(\sr_51_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_52_[6]_net_1 ));
    DFN1E1C0 \sr_21_[9]  (.D(\sr_20_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_21_[9]_net_1 ));
    DFN1E1C0 \sr_47_[12]  (.D(\sr_46_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_47_[12]_net_1 ));
    DFN1E1C0 \sr_22_[4]  (.D(\sr_21_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_22_[4]_net_1 ));
    DFN1E1C0 \sr_10_[1]  (.D(\sr_9_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_10_[1]_net_1 ));
    DFN1E1C0 \sr_5_[4]  (.D(\sr_4_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_5_[4]_net_1 ));
    DFN1E1C0 \sr_62_[6]  (.D(\sr_61_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_62_[6]_net_1 ));
    DFN1E1C0 \sr_58_[2]  (.D(\sr_57_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_58_[2]_net_1 ));
    DFN1E1C0 \sr_55_[0]  (.D(\sr_54_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_55_[0]_net_1 ));
    DFN1E1C0 \sr_27_[3]  (.D(\sr_26_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_27_[3]_net_1 ));
    DFN1E1C0 \sr_21_[1]  (.D(\sr_20_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_21_[1]_net_1 ));
    DFN1E1C0 \sr_37_[9]  (.D(\sr_36_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[9]_net_1 ));
    DFN1E1C0 \sr_48_[10]  (.D(\sr_47_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_48_[10]_net_1 ));
    DFN1E1C0 \sr_60_[5]  (.D(\sr_59_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_60_[5]_net_1 ));
    DFN1E1C0 \sr_30_[5]  (.D(\sr_29_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_30_[5]_net_1 ));
    DFN1E1C0 \sr_14_[4]  (.D(\sr_13_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_14_[4]_net_1 ));
    DFN1E1C0 \sr_24_[8]  (.D(\sr_23_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_24_[8]_net_1 ));
    DFN1E1C0 \sr_30_[4]  (.D(\sr_29_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_30_[4]_net_1 ));
    DFN1E1C0 \sr_37_[6]  (.D(\sr_36_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[6]_net_1 ));
    DFN1E1C0 \sr_42_[6]  (.D(\sr_41_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_42_[6]_net_1 ));
    DFN1E1C0 \sr_58_[4]  (.D(\sr_57_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_58_[4]_net_1 ));
    DFN1E1C0 \sr_57_[10]  (.D(\sr_56_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_5), .Q(\sr_57_[10]_net_1 ));
    DFN1E1C0 \sr_43_[7]  (.D(\sr_42_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_43_[7]_net_1 ));
    DFN1E1C0 \sr_44_[2]  (.D(\sr_43_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_44_[2]_net_1 ));
    DFN1E1C0 \sr_53_[7]  (.D(\sr_52_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_53_[7]_net_1 ));
    DFN1E1C0 \sr_59_[1]  (.D(\sr_58_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_59_[1]_net_1 ));
    DFN1E1C0 \sr_63__0[12]  (.D(\sr_62_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(sr_old_0_0));
    DFN1E1C0 \sr_27_[10]  (.D(\sr_26_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_27_[10]_net_1 ));
    DFN1E1C0 \sr_53_[8]  (.D(\sr_52_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_53_[8]_net_1 ));
    DFN1E1C0 \sr_16_[4]  (.D(\sr_15_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_16_[4]_net_1 ));
    DFN1E1C0 \sr_10_[11]  (.D(\sr_9_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_10_[11]_net_1 ));
    DFN1E1C0 \sr_26_[8]  (.D(\sr_25_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_26_[8]_net_1 ));
    DFN1E1C0 \sr_63_[7]  (.D(\sr_62_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[7]));
    DFN1E1C0 \sr_28_[7]  (.D(\sr_27_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_28_[7]_net_1 ));
    DFN1E1C0 \sr_63_[8]  (.D(\sr_62_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[8]));
    DFN1E1C0 \sr_24_[0]  (.D(\sr_23_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_24_[0]_net_1 ));
    DFN1E1C0 \sr_46_[2]  (.D(\sr_45_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_46_[2]_net_1 ));
    DFN1E1C0 \sr_13_[5]  (.D(\sr_12_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_13_[5]_net_1 ));
    DFN1E1C0 \sr_0_[2]  (.D(cur_error[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_21), .Q(sr_new[2]));
    DFN1E1C0 \sr_0_[8]  (.D(cur_error[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_21), .Q(sr_new[8]));
    DFN1E1C0 \sr_8_[3]  (.D(\sr_7_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_8_[3]_net_1 ));
    DFN1E1C0 \sr_42_[11]  (.D(\sr_41_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_42_[11]_net_1 ));
    DFN1E1C0 \sr_13_[3]  (.D(\sr_12_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_13_[3]_net_1 ));
    DFN1E1C0 \sr_54_[10]  (.D(\sr_53_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_54_[10]_net_1 ));
    DFN1E1C0 \sr_37_[11]  (.D(\sr_36_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_37_[11]_net_1 ));
    DFN1E1C0 \sr_19_[7]  (.D(\sr_18_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_19_[7]_net_1 ));
    DFN1E1C0 \sr_57_[1]  (.D(\sr_56_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_57_[1]_net_1 ));
    DFN1E1C0 \sr_44_[11]  (.D(\sr_43_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_44_[11]_net_1 ));
    DFN1E1C0 \sr_32_[10]  (.D(\sr_31_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_32_[10]_net_1 ));
    DFN1E1C0 \sr_26_[0]  (.D(\sr_25_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_26_[0]_net_1 ));
    DFN1E1C0 \sr_24_[10]  (.D(\sr_23_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_24_[10]_net_1 ));
    DFN1E1C0 \sr_12_[1]  (.D(\sr_11_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_12_[1]_net_1 ));
    DFN1E1C0 \sr_10_[4]  (.D(\sr_9_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_10_[4]_net_1 ));
    DFN1E1C0 \sr_63_[0]  (.D(\sr_62_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[0]));
    DFN1E1C0 \sr_20_[8]  (.D(\sr_19_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_20_[8]_net_1 ));
    DFN1E1C0 \sr_60_[12]  (.D(\sr_59_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_60_[12]_net_1 ));
    DFN1E1C0 \sr_6_[10]  (.D(\sr_5_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_6_[10]_net_1 ));
    DFN1E1C0 \sr_19_[6]  (.D(\sr_18_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_19_[6]_net_1 ));
    DFN1E1C0 \sr_62_[5]  (.D(\sr_61_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_62_[5]_net_1 ));
    DFN1E1C0 \sr_44_[8]  (.D(\sr_43_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_44_[8]_net_1 ));
    DFN1E1C0 \sr_49_[5]  (.D(\sr_48_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_49_[5]_net_1 ));
    DFN1E1C0 \sr_53_[0]  (.D(\sr_52_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_53_[0]_net_1 ));
    DFN1E1C0 \sr_1_[2]  (.D(sr_new[2]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable_30), .Q(sr_prev[2]));
    DFN1E1C0 \sr_40_[2]  (.D(\sr_39_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_40_[2]_net_1 ));
    DFN1E1C0 \sr_32_[5]  (.D(\sr_31_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_32_[5]_net_1 ));
    DFN1E1C0 \sr_1_[8]  (.D(sr_new[8]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable_31), .Q(sr_prev[8]));
    DFN1E1C0 \sr_18_[12]  (.D(\sr_17_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_18_[12]_net_1 ));
    DFN1E1C0 \sr_60_[10]  (.D(\sr_59_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_60_[10]_net_1 ));
    DFN1E1C0 \sr_32_[4]  (.D(\sr_31_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_32_[4]_net_1 ));
    DFN1E1C0 \sr_54_[3]  (.D(\sr_53_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_54_[3]_net_1 ));
    DFN1E1C0 \sr_29_[9]  (.D(\sr_28_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(\sr_29_[9]_net_1 ));
    DFN1E1C0 \sr_24_[2]  (.D(\sr_23_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_24_[2]_net_1 ));
    DFN1E1C0 \sr_18_[9]  (.D(\sr_17_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_18_[9]_net_1 ));
    DFN1E1C0 \sr_7_[9]  (.D(\sr_6_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_7_[9]_net_1 ));
    DFN1E1C0 \sr_63_[10]  (.D(\sr_62_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[10]));
    DFN1E1C0 \sr_24_[5]  (.D(\sr_23_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_24_[5]_net_1 ));
    DFN1E1C0 \sr_46_[8]  (.D(\sr_45_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_46_[8]_net_1 ));
    DFN1E1C0 \sr_59_[11]  (.D(\sr_58_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_59_[11]_net_1 ));
    DFN1E1C0 \sr_17_[7]  (.D(\sr_16_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_17_[7]_net_1 ));
    DFN1E1C0 \sr_14_[8]  (.D(\sr_13_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_14_[8]_net_1 ));
    DFN1E1C0 \sr_41_[3]  (.D(\sr_40_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_41_[3]_net_1 ));
    DFN1E1C0 \sr_20_[0]  (.D(\sr_19_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_20_[0]_net_1 ));
    DFN1E1C0 \sr_48_[0]  (.D(\sr_47_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_48_[0]_net_1 ));
    DFN1E1C0 \sr_29_[1]  (.D(\sr_28_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(\sr_29_[1]_net_1 ));
    DFN1E1C0 \sr_3_[10]  (.D(\sr_2_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_3_[10]_net_1 ));
    DFN1E1C0 \sr_29_[11]  (.D(\sr_28_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_29_[11]_net_1 ));
    DFN1E1C0 \sr_35_[1]  (.D(\sr_34_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_35_[1]_net_1 ));
    DFN1E1C0 \sr_17_[6]  (.D(\sr_16_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_17_[6]_net_1 ));
    DFN1E1C0 \sr_2_[3]  (.D(sr_prev[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_5), .Q(\sr_2_[3]_net_1 ));
    DFN1E1C0 \sr_56_[3]  (.D(\sr_55_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_56_[3]_net_1 ));
    DFN1E1C0 \sr_47_[5]  (.D(\sr_46_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_47_[5]_net_1 ));
    DFN1E1C0 \sr_35_[2]  (.D(\sr_34_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_35_[2]_net_1 ));
    DFN1E1C0 \sr_35_[12]  (.D(\sr_34_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_35_[12]_net_1 ));
    DFN1E1C0 \sr_26_[2]  (.D(\sr_25_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_26_[2]_net_1 ));
    DFN1E1C0 \sr_6_[2]  (.D(\sr_5_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_6_[2]_net_1 ));
    DFN1E1C0 \sr_6_[8]  (.D(\sr_5_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_6_[8]_net_1 ));
    DFN1E1C0 \sr_35_[7]  (.D(\sr_34_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_35_[7]_net_1 ));
    DFN1E1C0 \sr_26_[5]  (.D(\sr_25_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_26_[5]_net_1 ));
    DFN1E1C0 \sr_16_[8]  (.D(\sr_15_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_16_[8]_net_1 ));
    DFN1E1C0 \sr_52_[12]  (.D(\sr_51_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_52_[12]_net_1 ));
    DFN1E1C0 \sr_5_[2]  (.D(\sr_4_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_5_[2]_net_1 ));
    DFN1E1C0 \sr_5_[8]  (.D(\sr_4_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_5_[8]_net_1 ));
    DFN1E1C0 \sr_27_[9]  (.D(\sr_26_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_27_[9]_net_1 ));
    DFN1E1C0 \sr_18_[11]  (.D(\sr_17_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_18_[11]_net_1 ));
    DFN1E1C0 \sr_3_[9]  (.D(\sr_2_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_3_[9]_net_1 ));
    DFN1E1C0 \sr_2_[11]  (.D(sr_prev[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_14), .Q(\sr_2_[11]_net_1 ));
    DFN1E1C0 \sr_40_[8]  (.D(\sr_39_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_40_[8]_net_1 ));
    DFN1E1C0 \sr_22_[12]  (.D(\sr_21_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_22_[12]_net_1 ));
    DFN1E1C0 \sr_45_[9]  (.D(\sr_44_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_45_[9]_net_1 ));
    DFN1E1C0 \sr_2_[12]  (.D(sr_prev[12]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_14), .Q(\sr_2_[12]_net_1 ));
    DFN1E1C0 \sr_27_[1]  (.D(\sr_26_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_27_[1]_net_1 ));
    DFN1E1C0 \sr_0__1[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(sr_new_1_0));
    DFN1E1C0 \sr_9_[4]  (.D(\sr_8_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[4]_net_1 ));
    DFN1E1C0 \sr_12_[4]  (.D(\sr_11_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_12_[4]_net_1 ));
    DFN1E1C0 \sr_56_[11]  (.D(\sr_55_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_56_[11]_net_1 ));
    DFN1E1C0 \sr_22_[8]  (.D(\sr_21_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_22_[8]_net_1 ));
    DFN1E1C0 \sr_14_[2]  (.D(\sr_13_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_14_[2]_net_1 ));
    DFN1E1C0 \sr_46_[12]  (.D(\sr_45_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_46_[12]_net_1 ));
    DFN1E1C0 \sr_50_[3]  (.D(\sr_49_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_50_[3]_net_1 ));
    DFN1E1C0 \sr_20_[2]  (.D(\sr_19_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_20_[2]_net_1 ));
    DFN1E1C0 \sr_44_[12]  (.D(\sr_43_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_44_[12]_net_1 ));
    DFN1E1C0 \sr_26_[11]  (.D(\sr_25_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_26_[11]_net_1 ));
    DFN1E1C0 \sr_14_[0]  (.D(\sr_13_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_14_[0]_net_1 ));
    DFN1E1C0 \sr_34_[8]  (.D(\sr_33_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_34_[8]_net_1 ));
    DFN1E1C0 \sr_20_[5]  (.D(\sr_19_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_20_[5]_net_1 ));
    DFN1E1C0 \sr_10_[8]  (.D(\sr_9_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_10_[8]_net_1 ));
    DFN1E1C0 \sr_42_[2]  (.D(\sr_41_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_42_[2]_net_1 ));
    DFN1E1C0 \sr_55_[11]  (.D(\sr_54_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(\sr_55_[11]_net_1 ));
    DFN1E1C0 \sr_51_[9]  (.D(\sr_50_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_51_[9]_net_1 ));
    DFN1E1C0 \sr_54_[5]  (.D(\sr_53_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_54_[5]_net_1 ));
    DFN1E1C0 \sr_25_[11]  (.D(\sr_24_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_25_[11]_net_1 ));
    DFN1E1C0 \sr_21_[6]  (.D(\sr_20_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_21_[6]_net_1 ));
    DFN1E1C0 \sr_57_[12]  (.D(\sr_56_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_5), .Q(\sr_57_[12]_net_1 ));
    DFN1E1C0 \sr_16_[2]  (.D(\sr_15_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_16_[2]_net_1 ));
    DFN1E1C0 \sr_35_[0]  (.D(\sr_34_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_35_[0]_net_1 ));
    DFN1E1C0 \sr_16_[0]  (.D(\sr_15_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_16_[0]_net_1 ));
    DFN1E1C0 \sr_36_[8]  (.D(\sr_35_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_36_[8]_net_1 ));
    DFN1E1C0 \sr_27_[12]  (.D(\sr_26_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_27_[12]_net_1 ));
    DFN1E1C0 \sr_22_[0]  (.D(\sr_21_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_22_[0]_net_1 ));
    DFN1E1C0 \sr_0__0[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(sr_new_0_0));
    DFN1E1C0 \sr_13_[11]  (.D(\sr_12_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_13_[11]_net_1 ));
    DFN1E1C0 \sr_58_[10]  (.D(\sr_57_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_58_[10]_net_1 ));
    DFN1E1C0 \sr_7_[12]  (.D(\sr_6_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_7_[12]_net_1 ));
    DFN1E1C0 \sr_24_[3]  (.D(\sr_23_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_24_[3]_net_1 ));
    DFN1E1C0 \sr_34_[9]  (.D(\sr_33_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_34_[9]_net_1 ));
    DFN1E1C0 \sr_28_[10]  (.D(\sr_27_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_28_[10]_net_1 ));
    DFN1E1C0 \sr_56_[5]  (.D(\sr_55_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_56_[5]_net_1 ));
    DFN1E1C0 \sr_7_[10]  (.D(\sr_6_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_7_[10]_net_1 ));
    DFN1E1C0 \sr_33_[1]  (.D(\sr_32_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_33_[1]_net_1 ));
    DFN1E1C0 \sr_33_[2]  (.D(\sr_32_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_33_[2]_net_1 ));
    DFN1E1C0 \sr_48_[7]  (.D(\sr_47_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_48_[7]_net_1 ));
    DFN1E1C0 \sr_58_[7]  (.D(\sr_57_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_58_[7]_net_1 ));
    DFN1E1C0 \sr_34_[6]  (.D(\sr_33_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_34_[6]_net_1 ));
    DFN1E1C0 \sr_33_[7]  (.D(\sr_32_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_33_[7]_net_1 ));
    DFN1E1C0 \sr_10_[2]  (.D(\sr_9_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_10_[2]_net_1 ));
    DFN1E1C0 \sr_26_[3]  (.D(\sr_25_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_26_[3]_net_1 ));
    DFN1E1C0 \sr_36_[9]  (.D(\sr_35_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_36_[9]_net_1 ));
    DFN1E1C0 \sr_58_[8]  (.D(\sr_57_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_58_[8]_net_1 ));
    DFN1E1C0 \sr_42_[8]  (.D(\sr_41_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_42_[8]_net_1 ));
    DFN1E1C0 \sr_49_[3]  (.D(\sr_48_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_49_[3]_net_1 ));
    DFN1E1C0 \sr_10_[0]  (.D(\sr_9_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_10_[0]_net_1 ));
    DFN1E1C0 \sr_30_[8]  (.D(\sr_29_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_30_[8]_net_1 ));
    DFN1E1C0 \sr_35_[10]  (.D(\sr_34_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_35_[10]_net_1 ));
    DFN1E1C0 \sr_8_[4]  (.D(\sr_7_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_8_[4]_net_1 ));
    DFN1E1C0 \sr_43_[12]  (.D(\sr_42_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_43_[12]_net_1 ));
    DFN1E1C0 \sr_0_[9]  (.D(cur_error[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_21), .Q(sr_new[9]));
    DFN1E1C0 \sr_43_[9]  (.D(\sr_42_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_43_[9]_net_1 ));
    DFN1E1C0 \sr_50_[5]  (.D(\sr_49_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_50_[5]_net_1 ));
    DFN1E1C0 \sr_52_[3]  (.D(\sr_51_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_52_[3]_net_1 ));
    DFN1E1C0 \sr_22_[2]  (.D(\sr_21_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_22_[2]_net_1 ));
    DFN1E1C0 \sr_18_[5]  (.D(\sr_17_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_18_[5]_net_1 ));
    DFN1E1C0 \sr_7_[0]  (.D(\sr_6_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_7_[0]_net_1 ));
    DFN1E1C0 \sr_36_[6]  (.D(\sr_35_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_36_[6]_net_1 ));
    DFN1E1C0 \sr_60_[11]  (.D(\sr_59_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_60_[11]_net_1 ));
    DFN1E1C0 \sr_45_[4]  (.D(\sr_44_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_45_[4]_net_1 ));
    DFN1E1C0 \sr_22_[5]  (.D(\sr_21_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_22_[5]_net_1 ));
    DFN1E1C0 \sr_35_[3]  (.D(\sr_34_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_35_[3]_net_1 ));
    DFN1E1C0 \sr_7_[6]  (.D(\sr_6_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_7_[6]_net_1 ));
    DFN1E1C0 \sr_12_[8]  (.D(\sr_11_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_12_[8]_net_1 ));
    DFN1E1C0 \sr_55_[6]  (.D(\sr_54_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_55_[6]_net_1 ));
    DFN1E1C0 \sr_52_[11]  (.D(\sr_51_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_52_[11]_net_1 ));
    DFN1E1C0 \sr_18_[3]  (.D(\sr_17_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_18_[3]_net_1 ));
    DFN1E1C0 \sr_36_[10]  (.D(\sr_35_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_36_[10]_net_1 ));
    DFN1E1C0 \sr_25_[4]  (.D(\sr_24_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_25_[4]_net_1 ));
    DFN1E1C0 \sr_22_[11]  (.D(\sr_21_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_22_[11]_net_1 ));
    DFN1E1C0 \sr_20_[3]  (.D(\sr_19_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_20_[3]_net_1 ));
    DFN1E1C0 \sr_30_[9]  (.D(\sr_29_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_30_[9]_net_1 ));
    DFN1E1C0 \sr_47_[3]  (.D(\sr_46_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_47_[3]_net_1 ));
    DFN1E1C0 \sr_54_[11]  (.D(\sr_53_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_54_[11]_net_1 ));
    DFN1E1C0 \sr_4_[7]  (.D(\sr_3_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_4_[7]_net_1 ));
    DFN1E1C0 \sr_31_[12]  (.D(\sr_30_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_31_[12]_net_1 ));
    DFN1E1C0 \sr_54_[1]  (.D(\sr_53_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_54_[1]_net_1 ));
    DFN1E1C0 \sr_24_[11]  (.D(\sr_23_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_24_[11]_net_1 ));
    DFN1E1C0 \sr_1_[9]  (.D(sr_new[9]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable_31), .Q(sr_prev[9]));
    DFN1E1C0 \sr_58_[0]  (.D(\sr_57_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_58_[0]_net_1 ));
    DFN1E1C0 \sr_33_[0]  (.D(\sr_32_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_33_[0]_net_1 ));
    DFN1E1C0 \sr_41_[1]  (.D(\sr_40_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_41_[1]_net_1 ));
    DFN1E1C0 \sr_30_[6]  (.D(\sr_29_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_30_[6]_net_1 ));
    DFN1E1C0 \sr_7_[1]  (.D(\sr_6_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_7_[1]_net_1 ));
    DFN1E1C0 \sr_3_[0]  (.D(\sr_2_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_3_[0]_net_1 ));
    DFN1E1C0 \sr_45_[6]  (.D(\sr_44_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_45_[6]_net_1 ));
    DFN1E1C0 \sr_3_[6]  (.D(\sr_2_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_3_[6]_net_1 ));
    DFN1E1C0 \sr_59_[9]  (.D(\sr_58_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_59_[9]_net_1 ));
    DFN1E1C0 \sr_2_[4]  (.D(sr_prev[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_5), .Q(\sr_2_[4]_net_1 ));
    DFN1E1C0 \sr_56_[1]  (.D(\sr_55_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_56_[1]_net_1 ));
    DFN1E1C0 \sr_29_[6]  (.D(\sr_28_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(\sr_29_[6]_net_1 ));
    DFN1E1C0 \sr_9_[2]  (.D(\sr_8_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[2]_net_1 ));
    DFN1E1C0 \sr_9_[8]  (.D(\sr_8_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[8]_net_1 ));
    DFN1E1C0 \sr_17_[11]  (.D(\sr_16_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_17_[11]_net_1 ));
    DFN1E1C0 \sr_12_[2]  (.D(\sr_11_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_12_[2]_net_1 ));
    DFN1E1C0 \sr_12_[10]  (.D(\sr_11_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_12_[10]_net_1 ));
    DFN1E1C0 \sr_12_[0]  (.D(\sr_11_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_12_[0]_net_1 ));
    DFN1E1C0 \sr_32_[8]  (.D(\sr_31_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_32_[8]_net_1 ));
    DFN1E1C0 \sr_14_[7]  (.D(\sr_13_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_14_[7]_net_1 ));
    DFN1E1C0 \sr_6_[9]  (.D(\sr_5_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_6_[9]_net_1 ));
    DFN1E1C0 \sr_31_[10]  (.D(\sr_30_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_31_[10]_net_1 ));
    DFN1E1C0 \sr_31_[11]  (.D(\sr_30_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_31_[11]_net_1 ));
    DFN1E1C0 \sr_14_[6]  (.D(\sr_13_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_14_[6]_net_1 ));
    DFN1E1C0 \sr_5_[10]  (.D(\sr_4_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_5_[10]_net_1 ));
    DFN1E1C0 \sr_5_[9]  (.D(\sr_4_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_5_[9]_net_1 ));
    DFN1E1C0 \sr_52_[5]  (.D(\sr_51_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_52_[5]_net_1 ));
    DFN1E1C0 \sr_3_[1]  (.D(\sr_2_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_3_[1]_net_1 ));
    DFN1E1C0 \sr_44_[5]  (.D(\sr_43_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_44_[5]_net_1 ));
    DFN1E1C0 \sr_57_[9]  (.D(\sr_56_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_57_[9]_net_1 ));
    DFN1E1C0 \sr_50_[1]  (.D(\sr_49_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_50_[1]_net_1 ));
    DFN1E1C0 \sr_16_[7]  (.D(\sr_15_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_16_[7]_net_1 ));
    DFN1E1C0 \sr_51_[2]  (.D(\sr_50_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_51_[2]_net_1 ));
    DFN1E1C0 \sr_27_[6]  (.D(\sr_26_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_27_[6]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1C0 \sr_43_[4]  (.D(\sr_42_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_43_[4]_net_1 ));
    DFN1E1C0 \sr_24_[9]  (.D(\sr_23_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_24_[9]_net_1 ));
    DFN1E1C0 \sr_22_[3]  (.D(\sr_21_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_22_[3]_net_1 ));
    DFN1E1C0 \sr_33_[3]  (.D(\sr_32_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_33_[3]_net_1 ));
    DFN1E1C0 \sr_32_[9]  (.D(\sr_31_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_32_[9]_net_1 ));
    DFN1E1C0 \sr_15_[1]  (.D(\sr_14_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_5), .Q(\sr_15_[1]_net_1 ));
    DFN1E1C0 \sr_53_[6]  (.D(\sr_52_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_53_[6]_net_1 ));
    DFN1E1C0 \sr_60_[1]  (.D(\sr_59_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_60_[1]_net_1 ));
    DFN1E1C0 \sr_16_[6]  (.D(\sr_15_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_16_[6]_net_1 ));
    DFN1E1C0 \sr_61_[2]  (.D(\sr_60_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_61_[2]_net_1 ));
    DFN1E1C0 \sr_23_[4]  (.D(\sr_22_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_23_[4]_net_1 ));
    DFN1E1C0 \sr_46_[5]  (.D(\sr_45_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_46_[5]_net_1 ));
    DFN1E1C0 \sr_24_[1]  (.D(\sr_23_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_24_[1]_net_1 ));
    DFN1E1C0 \sr_63_[6]  (.D(\sr_62_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[6]));
    DFN1E1C0 \sr_49_[12]  (.D(\sr_48_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_49_[12]_net_1 ));
    DFN1E1C0 \sr_56_[12]  (.D(\sr_55_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_56_[12]_net_1 ));
    DFN1E1C0 \sr_54_[12]  (.D(\sr_53_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_54_[12]_net_1 ));
    DFN1E1C0 \sr_35_[5]  (.D(\sr_34_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_35_[5]_net_1 ));
    DFN1E1C0 \sr_15_[12]  (.D(\sr_14_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_15_[12]_net_1 ));
    DFN1E1C0 \sr_32_[6]  (.D(\sr_31_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_32_[6]_net_1 ));
    DFN1E1C0 \sr_26_[12]  (.D(\sr_25_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_26_[12]_net_1 ));
    DFN1E1C0 \sr_35_[4]  (.D(\sr_34_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_35_[4]_net_1 ));
    DFN1E1C0 \sr_26_[9]  (.D(\sr_25_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_26_[9]_net_1 ));
    DFN1E1C0 \sr_24_[12]  (.D(\sr_23_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_24_[12]_net_1 ));
    DFN1E1C0 \sr_51_[4]  (.D(\sr_50_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_51_[4]_net_1 ));
    DFN1E1C0 \sr_10_[7]  (.D(\sr_9_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_10_[7]_net_1 ));
    DFN1E1C0 \sr_8_[2]  (.D(\sr_7_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_8_[2]_net_1 ));
    DFN1E1C0 \sr_40_[12]  (.D(\sr_39_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_40_[12]_net_1 ));
    DFN1E1C0 \sr_8_[8]  (.D(\sr_7_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_8_[8]_net_1 ));
    DFN1E1C0 \sr_26_[1]  (.D(\sr_25_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_26_[1]_net_1 ));
    DFN1E1C0 \sr_61_[4]  (.D(\sr_60_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_61_[4]_net_1 ));
    DFN1E1C0 \sr_0_[0]  (.D(cur_error[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_20), .Q(sr_new[0]));
    DFN1E1C0 \sr_43_[6]  (.D(\sr_42_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_43_[6]_net_1 ));
    DFN1E1C0 \sr_10_[6]  (.D(\sr_9_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_10_[6]_net_1 ));
    DFN1E1C0 \sr_21_[7]  (.D(\sr_20_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_21_[7]_net_1 ));
    DFN1E1C0 \sr_0_[6]  (.D(cur_error[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_21), .Q(sr_new[6]));
    DFN1E1C0 \sr_40_[5]  (.D(\sr_39_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_40_[5]_net_1 ));
    DFN1E1C0 \sr_40_[10]  (.D(\sr_39_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_40_[10]_net_1 ));
    DFN1E1C0 \sr_43_[10]  (.D(\sr_42_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_43_[10]_net_1 ));
    DFN1E1C0 \sr_38_[1]  (.D(\sr_37_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[1]_net_1 ));
    DFN1E1C0 \sr_49_[1]  (.D(\sr_48_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_49_[1]_net_1 ));
    DFN1E1C0 \sr_63_[11]  (.D(\sr_62_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[11]));
    DFN1E1C0 \sr_20_[9]  (.D(\sr_19_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_20_[9]_net_1 ));
    DFN1E1C0 \sr_38_[2]  (.D(\sr_37_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[2]_net_1 ));
    DFN1E1C0 \sr_38_[7]  (.D(\sr_37_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[7]_net_1 ));
    DFN1E1C0 \sr_52_[1]  (.D(\sr_51_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_52_[1]_net_1 ));
    DFN1E1C0 \sr_20_[1]  (.D(\sr_19_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_20_[1]_net_1 ));
    DFN1E1C0 \sr_1_[0]  (.D(sr_new[0]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable_30), .Q(sr_prev[0]));
    DFN1E1C0 \sr_61_[9]  (.D(\sr_60_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_61_[9]_net_1 ));
    DFN1E1C0 \sr_0_[1]  (.D(cur_error[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_21), .Q(sr_new[1]));
    DFN1E1C0 \sr_15_[4]  (.D(\sr_14_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_5), .Q(\sr_15_[4]_net_1 ));
    DFN1E1C0 \sr_1_[6]  (.D(sr_new[6]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable_30), .Q(sr_prev[6]));
    DFN1E1C0 \sr_62_[1]  (.D(\sr_61_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_62_[1]_net_1 ));
    DFN1E1C0 \sr_25_[8]  (.D(\sr_24_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_25_[8]_net_1 ));
    DFN1E1C0 \sr_48_[9]  (.D(\sr_47_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_48_[9]_net_1 ));
    DFN1E1C0 \sr_1_[11]  (.D(sr_new[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_27), .Q(sr_prev[11]));
    DFN1E1C0 \sr_49_[10]  (.D(\sr_48_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_49_[10]_net_1 ));
    DFN1E1C0 \sr_53_[12]  (.D(\sr_52_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_53_[12]_net_1 ));
    DFN1E1C0 \sr_13_[1]  (.D(\sr_12_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_13_[1]_net_1 ));
    DFN1E1C0 \sr_7_[5]  (.D(\sr_6_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_7_[5]_net_1 ));
    DFN1E1C0 \sr_5_[12]  (.D(\sr_4_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_5_[12]_net_1 ));
    DFN1E1C0 \sr_47_[1]  (.D(\sr_46_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_47_[1]_net_1 ));
    DFN1E1C0 \sr_23_[12]  (.D(\sr_22_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_23_[12]_net_1 ));
    DFN1E1C0 \sr_63_[5]  (.D(\sr_62_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[5]));
    DFN1E1C0 \sr_45_[2]  (.D(\sr_44_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_45_[2]_net_1 ));
    DFN1E1C0 \sr_2_[2]  (.D(sr_prev[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_5), .Q(\sr_2_[2]_net_1 ));
    DFN1E1C0 \sr_2_[8]  (.D(sr_prev[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_5), .Q(\sr_2_[8]_net_1 ));
    DFN1E1C0 \sr_11_[9]  (.D(\sr_10_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_11_[9]_net_1 ));
    DFN1E1C0 \sr_33_[5]  (.D(\sr_32_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_33_[5]_net_1 ));
    DFN1E1C0 \sr_59_[2]  (.D(\sr_58_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_59_[2]_net_1 ));
    DFN1E1C0 \sr_12_[7]  (.D(\sr_11_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_12_[7]_net_1 ));
    DFN1E1C0 \sr_6_[0]  (.D(\sr_5_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_6_[0]_net_1 ));
    DFN1E1C0 \sr_41_[0]  (.D(\sr_40_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_41_[0]_net_1 ));
    DFN1E1C0 \sr_1_[1]  (.D(sr_new[1]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable_30), .Q(sr_prev[1]));
    DFN1E1C0 \sr_33_[4]  (.D(\sr_32_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_33_[4]_net_1 ));
    DFN1E1C0 \sr_9_[12]  (.D(\sr_8_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_9_[12]_net_1 ));
    DFN1E1C0 \sr_25_[0]  (.D(\sr_24_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_25_[0]_net_1 ));
    DFN1E1C0 \sr_6_[6]  (.D(\sr_5_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_6_[6]_net_1 ));
    DFN1E1C0 \sr_15_[10]  (.D(\sr_14_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_15_[10]_net_1 ));
    DFN1E1C0 \sr_12_[6]  (.D(\sr_11_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_12_[6]_net_1 ));
    DFN1E1C0 \sr_61_[3]  (.D(\sr_60_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_61_[3]_net_1 ));
    DFN1E1C0 \sr_5_[0]  (.D(\sr_4_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_5_[0]_net_1 ));
    DFN1E1C0 \sr_44_[3]  (.D(\sr_43_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_44_[3]_net_1 ));
    DFN1E1C0 \sr_38_[0]  (.D(\sr_37_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[0]_net_1 ));
    DFN1E1C0 \sr_42_[5]  (.D(\sr_41_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_42_[5]_net_1 ));
    DFN1E1C0 \sr_5_[6]  (.D(\sr_4_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_5_[6]_net_1 ));
    DFN1E1C0 \sr_3_[5]  (.D(\sr_2_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_3_[5]_net_1 ));
    DFN1E1C0 \sr_4_[3]  (.D(\sr_3_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_4_[3]_net_1 ));
    DFN1E1C0 \sr_9_[9]  (.D(\sr_8_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[9]_net_1 ));
    DFN1E1C0 \sr_37_[10]  (.D(\sr_36_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_37_[10]_net_1 ));
    DFN1E1C0 \sr_22_[9]  (.D(\sr_21_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_22_[9]_net_1 ));
    DFN1E1C0 \sr_59_[4]  (.D(\sr_58_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_59_[4]_net_1 ));
    DFN1E1C0 \sr_16_[10]  (.D(\sr_15_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_16_[10]_net_1 ));
    DFN1E1C0 \sr_57_[2]  (.D(\sr_56_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_57_[2]_net_1 ));
    DFN1E1C0 \sr_46_[3]  (.D(\sr_45_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_46_[3]_net_1 ));
    DFN1E1C0 \sr_6_[1]  (.D(\sr_5_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_6_[1]_net_1 ));
    DFN1E1C0 \sr_45_[8]  (.D(\sr_44_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_45_[8]_net_1 ));
    DFN1E1C0 \sr_22_[1]  (.D(\sr_21_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_22_[1]_net_1 ));
    DFN1E1C0 \sr_29_[7]  (.D(\sr_28_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(\sr_29_[7]_net_1 ));
    DFN1E1C0 \sr_11_[12]  (.D(\sr_10_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_11_[12]_net_1 ));
    DFN1E1C0 \sr_5_[1]  (.D(\sr_4_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_5_[1]_net_1 ));
    DFN1E1C0 \sr_4_[10]  (.D(\sr_3_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_4_[10]_net_1 ));
    DFN1E1C0 \sr_55_[3]  (.D(\sr_54_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_55_[3]_net_1 ));
    DFN1E1C0 \sr_25_[2]  (.D(\sr_24_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_25_[2]_net_1 ));
    DFN1E1C0 \sr_13_[4]  (.D(\sr_12_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_13_[4]_net_1 ));
    DFN1E1C0 \sr_62_[10]  (.D(\sr_61_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_62_[10]_net_1 ));
    DFN1E1C0 \sr_23_[8]  (.D(\sr_22_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_23_[8]_net_1 ));
    DFN1E1C0 \sr_25_[5]  (.D(\sr_24_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_25_[5]_net_1 ));
    DFN1E1C0 \sr_15_[8]  (.D(\sr_14_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_15_[8]_net_1 ));
    DFN1E1C0 \sr_34_[10]  (.D(\sr_33_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_34_[10]_net_1 ));
    DFN1E1C0 \sr_57_[4]  (.D(\sr_56_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_57_[4]_net_1 ));
    DFN1E1C0 \sr_40_[3]  (.D(\sr_39_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_40_[3]_net_1 ));
    DFN1E1C0 \sr_48_[4]  (.D(\sr_47_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_48_[4]_net_1 ));
    DFN1E1C0 \sr_38_[3]  (.D(\sr_37_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[3]_net_1 ));
    DFN1E1C0 \sr_43_[2]  (.D(\sr_42_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_43_[2]_net_1 ));
    DFN1E1C0 \sr_58_[6]  (.D(\sr_57_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_58_[6]_net_1 ));
    DFN1E1C0 \sr_54_[9]  (.D(\sr_53_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_54_[9]_net_1 ));
    DFN1E1C0 \sr_28_[4]  (.D(\sr_27_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_28_[4]_net_1 ));
    DFN1E1C0 \sr_27_[7]  (.D(\sr_26_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_27_[7]_net_1 ));
    DFN1E1C0 \sr_24_[6]  (.D(\sr_23_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_24_[6]_net_1 ));
    DFN1E1C0 \sr_40_[11]  (.D(\sr_39_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_40_[11]_net_1 ));
    DFN1E1C0 \sr_11_[10]  (.D(\sr_10_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_11_[10]_net_1 ));
    DFN1E1C0 \sr_23_[0]  (.D(\sr_22_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_23_[0]_net_1 ));
    DFN1E1C0 \sr_11_[11]  (.D(\sr_10_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_11_[11]_net_1 ));
    DFN1E1C0 \sr_59_[12]  (.D(\sr_58_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_59_[12]_net_1 ));
    DFN1E1C0 \sr_8_[9]  (.D(\sr_7_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_8_[9]_net_1 ));
    DFN1E1C0 \sr_1_[10]  (.D(sr_new[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_27), .Q(sr_prev[10]));
    DFN1E1C0 \sr_41_[7]  (.D(\sr_40_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_41_[7]_net_1 ));
    DFN1E1C0 \sr_29_[12]  (.D(\sr_28_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_29_[12]_net_1 ));
    DFN1E1C0 \sr_19_[9]  (.D(\sr_18_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_19_[9]_net_1 ));
    DFN1E1C0 \sr_56_[9]  (.D(\sr_55_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_56_[9]_net_1 ));
    DFN1E1C0 \sr_51_[7]  (.D(\sr_50_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_51_[7]_net_1 ));
    DFN1E1C0 \sr_39_[11]  (.D(\sr_38_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_39_[11]_net_1 ));
    DFN1E1C0 \sr_26_[6]  (.D(\sr_25_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_26_[6]_net_1 ));
    DFN1E1C0 \sr_51_[8]  (.D(\sr_50_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_51_[8]_net_1 ));
    DFN1E1C0 \sr_50_[12]  (.D(\sr_49_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_50_[12]_net_1 ));
    DFN1E1C0 \sr_49_[0]  (.D(\sr_48_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_49_[0]_net_1 ));
    DFN1E1C0 \sr_0_[5]  (.D(cur_error[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_21), .Q(sr_new[5]));
    DFN1E1C0 \sr_15_[2]  (.D(\sr_14_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_5), .Q(\sr_15_[2]_net_1 ));
    DFN1E1C0 \sr_61_[7]  (.D(\sr_60_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_61_[7]_net_1 ));
    DFN1E1C0 \sr_48_[6]  (.D(\sr_47_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_48_[6]_net_1 ));
    DFN1E1C0 \sr_15_[0]  (.D(\sr_14_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_5), .Q(\sr_15_[0]_net_1 ));
    DFN1E1C0 \sr_35_[8]  (.D(\sr_34_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_35_[8]_net_1 ));
    DFN1E1C0 \sr_61_[8]  (.D(\sr_60_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_61_[8]_net_1 ));
    DFN1E1C0 \sr_20_[12]  (.D(\sr_19_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_20_[12]_net_1 ));
    DFN1E1C0 \sr_43_[8]  (.D(\sr_42_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_43_[8]_net_1 ));
    DFN1E1C0 \sr_11_[5]  (.D(\sr_10_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_11_[5]_net_1 ));
    DFN1E1C0 \sr_50_[10]  (.D(\sr_49_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_50_[10]_net_1 ));
    DFN1E1C0 \sr_55_[5]  (.D(\sr_54_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_55_[5]_net_1 ));
    DFN1E1C0 \sr_53_[10]  (.D(\sr_52_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_53_[10]_net_1 ));
    DFN1E1C0 \sr_48_[12]  (.D(\sr_47_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_48_[12]_net_1 ));
    DFN1E1C0 \sr_32_[12]  (.D(\sr_31_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_32_[12]_net_1 ));
    DFN1E1C0 \sr_11_[3]  (.D(\sr_10_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_11_[3]_net_1 ));
    DFN1E1C0 \sr_0_[11]  (.D(cur_error[11]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable_5), .Q(sr_new[11]));
    DFN1E1C0 \sr_20_[10]  (.D(\sr_19_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_20_[10]_net_1 ));
    DFN1E1C0 \sr_50_[9]  (.D(\sr_49_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_50_[9]_net_1 ));
    DFN1E1C0 \sr_17_[9]  (.D(\sr_16_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_17_[9]_net_1 ));
    DFN1E1C0 \sr_23_[10]  (.D(\sr_22_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_23_[10]_net_1 ));
    DFN1E1C0 \sr_20_[6]  (.D(\sr_19_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_20_[6]_net_1 ));
    DFN1E1C0 \sr_53_[3]  (.D(\sr_52_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_53_[3]_net_1 ));
    DFN1E1C0 \sr_23_[2]  (.D(\sr_22_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_23_[2]_net_1 ));
    DFN1E1C0 \sr_1_[5]  (.D(sr_new[5]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable_30), .Q(sr_prev[5]));
    DFN1E1C0 \sr_61_[0]  (.D(\sr_60_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_61_[0]_net_1 ));
    DFN1E1C0 \sr_47_[0]  (.D(\sr_46_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_47_[0]_net_1 ));
    DFN1E1C0 \sr_23_[5]  (.D(\sr_22_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_23_[5]_net_1 ));
    DFN1E1C0 \sr_42_[3]  (.D(\sr_41_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_42_[3]_net_1 ));
    DFN1E1C0 \sr_25_[3]  (.D(\sr_24_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_25_[3]_net_1 ));
    DFN1E1C0 \sr_35_[9]  (.D(\sr_34_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_35_[9]_net_1 ));
    DFN1E1C0 \sr_13_[8]  (.D(\sr_12_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_13_[8]_net_1 ));
    DFN1E1C0 \sr_36_[11]  (.D(\sr_35_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_36_[11]_net_1 ));
    DFN1E1C0 \sr_51_[0]  (.D(\sr_50_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_51_[0]_net_1 ));
    DFN1E1C0 \sr_18_[1]  (.D(\sr_17_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_18_[1]_net_1 ));
    DFN1E1C0 \sr_2_[9]  (.D(sr_prev[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_5), .Q(\sr_2_[9]_net_1 ));
    DFN1E1C0 \sr_9_[0]  (.D(\sr_8_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[0]_net_1 ));
    DFN1E1C0 \sr_59_[10]  (.D(\sr_58_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_59_[10]_net_1 ));
    DFN1E1C0 \sr_35_[11]  (.D(\sr_34_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_35_[11]_net_1 ));
    DFN1E1C0 \sr_35_[6]  (.D(\sr_34_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_35_[6]_net_1 ));
    DFN1E1C0 \sr_9_[6]  (.D(\sr_8_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[6]_net_1 ));
    DFN1E1C0 \sr_29_[10]  (.D(\sr_28_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_29_[10]_net_1 ));
    DFN1E1C0 \sr_44_[1]  (.D(\sr_43_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_44_[1]_net_1 ));
    DFN1E1C0 \sr_38_[5]  (.D(\sr_37_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[5]_net_1 ));
    DFN1E1C0 \sr_37_[12]  (.D(\sr_36_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_37_[12]_net_1 ));
    DFN1E1C0 \sr_6_[5]  (.D(\sr_5_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_6_[5]_net_1 ));
    DFN1E1C0 \sr_48_[11]  (.D(\sr_47_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_48_[11]_net_1 ));
    DFN1E1C0 \sr_38_[4]  (.D(\sr_37_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[4]_net_1 ));
    DFN1E1C0 \sr_4_[4]  (.D(\sr_3_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_4_[4]_net_1 ));
    DFN1E1C0 \sr_38_[10]  (.D(\sr_37_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[10]_net_1 ));
    DFN1E1C0 \sr_5_[5]  (.D(\sr_4_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_5_[5]_net_1 ));
    DFN1E1C0 \sr_13_[2]  (.D(\sr_12_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_13_[2]_net_1 ));
    DFN1E1C0 \sr_46_[1]  (.D(\sr_45_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_46_[1]_net_1 ));
    DFN1E1C0 \sr_9_[1]  (.D(\sr_8_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[1]_net_1 ));
    DFN1E1C0 \sr_13_[0]  (.D(\sr_12_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_13_[0]_net_1 ));
    DFN1E1C0 \sr_33_[8]  (.D(\sr_32_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_33_[8]_net_1 ));
    DFN1E1C0 \sr_49_[7]  (.D(\sr_48_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_49_[7]_net_1 ));
    DFN1E1C0 \sr_59_[7]  (.D(\sr_58_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_59_[7]_net_1 ));
    DFN1E1C0 \sr_52_[9]  (.D(\sr_51_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_52_[9]_net_1 ));
    DFN1E1C0 \sr_59_[8]  (.D(\sr_58_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_59_[8]_net_1 ));
    DFN1E1C0 \sr_53_[5]  (.D(\sr_52_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_53_[5]_net_1 ));
    DFN1E1C0 \sr_22_[6]  (.D(\sr_21_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_22_[6]_net_1 ));
    DFN1E1C0 \sr_55_[1]  (.D(\sr_54_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_55_[1]_net_1 ));
    DFN1E1C0 \sr_54_[2]  (.D(\sr_53_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_54_[2]_net_1 ));
    DFN1E1C0 \sr_43_[11]  (.D(\sr_42_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_43_[11]_net_1 ));
    DFN1E1C0 \sr_8_[0]  (.D(\sr_7_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_8_[0]_net_1 ));
    DFN1E1C0 \sr_23_[3]  (.D(\sr_22_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_23_[3]_net_1 ));
    DFN1E1C0 \sr_40_[1]  (.D(\sr_39_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_40_[1]_net_1 ));
    DFN1E1C0 \sr_33_[9]  (.D(\sr_32_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_33_[9]_net_1 ));
    DFN1E1C0 \sr_19_[5]  (.D(\sr_18_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_19_[5]_net_1 ));
    DFN1E1C0 \sr_18_[4]  (.D(\sr_17_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_18_[4]_net_1 ));
    DFN1E1C0 \sr_28_[8]  (.D(\sr_27_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_28_[8]_net_1 ));
    DFN1E1C0 \sr_8_[6]  (.D(\sr_7_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_8_[6]_net_1 ));
    DFN1E1C0 \sr_32_[11]  (.D(\sr_31_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_32_[11]_net_1 ));
    DFN1E1C0 \sr_61_[12]  (.D(\sr_60_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_61_[12]_net_1 ));
    DFN1E1C0 \sr_19_[3]  (.D(\sr_18_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_19_[3]_net_1 ));
    DFN1E1C0 \sr_8_[11]  (.D(\sr_7_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_8_[11]_net_1 ));
    DFN1E1C0 \sr_47_[7]  (.D(\sr_46_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_47_[7]_net_1 ));
    DFN1E1C0 \sr_57_[7]  (.D(\sr_56_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_57_[7]_net_1 ));
    DFN1E1C0 \sr_56_[2]  (.D(\sr_55_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_56_[2]_net_1 ));
    DFN1E1C0 \sr_17_[10]  (.D(\sr_16_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_17_[10]_net_1 ));
    DFN1E1C0 \sr_57_[8]  (.D(\sr_56_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_57_[8]_net_1 ));
    DFN1E1C0 \sr_48_[2]  (.D(\sr_47_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_48_[2]_net_1 ));
    DFN1E1C0 \sr_15_[7]  (.D(\sr_14_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_5), .Q(\sr_15_[7]_net_1 ));
    DFN1E1C0 \sr_34_[11]  (.D(\sr_33_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_34_[11]_net_1 ));
    DFN1E1C0 \sr_33_[6]  (.D(\sr_32_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_33_[6]_net_1 ));
    DFN1E1C0 \sr_54_[4]  (.D(\sr_53_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_54_[4]_net_1 ));
    DFN1E1C0 \sr_15_[6]  (.D(\sr_14_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_5), .Q(\sr_15_[6]_net_1 ));
    DFN1E1C0 \sr_59_[0]  (.D(\sr_58_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_59_[0]_net_1 ));
    DFN1E1C0 \sr_50_[11]  (.D(\sr_49_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_50_[11]_net_1 ));
    DFN1E1C0 \sr_45_[5]  (.D(\sr_44_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_45_[5]_net_1 ));
    DFN1E1C0 \sr_8_[1]  (.D(\sr_7_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_8_[1]_net_1 ));
    DFN1E1C0 \sr_31_[1]  (.D(\sr_30_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_31_[1]_net_1 ));
    DFN1E1C0 \sr_28_[0]  (.D(\sr_27_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_28_[0]_net_1 ));
    DFN1E1C0 \sr_17_[5]  (.D(\sr_16_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_17_[5]_net_1 ));
    DFN1E1C0 \sr_24_[7]  (.D(\sr_23_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_24_[7]_net_1 ));
    DFN1E1C0 \sr_20_[11]  (.D(\sr_19_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_20_[11]_net_1 ));
    DFN1E1C0 \sr_31_[2]  (.D(\sr_30_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_31_[2]_net_1 ));
    DFN1E1C0 \sr_17_[3]  (.D(\sr_16_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_17_[3]_net_1 ));
    DFN1E1C0 \sr_56_[4]  (.D(\sr_55_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_56_[4]_net_1 ));
    DFN1E1C0 \sr_31_[7]  (.D(\sr_30_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_31_[7]_net_1 ));
    DFN1E1C0 \sr_25_[9]  (.D(\sr_24_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_25_[9]_net_1 ));
    DFN1E1C0 \sr_61_[10]  (.D(\sr_60_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_61_[10]_net_1 ));
    DFN1E1C0 \sr_50_[2]  (.D(\sr_49_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_50_[2]_net_1 ));
    DFN1E1C0 \sr_14_[10]  (.D(\sr_13_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_14_[10]_net_1 ));
    DFN1E1C0 \sr_61_[11]  (.D(\sr_60_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_61_[11]_net_1 ));
    DFN1E1C0 \sr_25_[1]  (.D(\sr_24_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_25_[1]_net_1 ));
    DFN1E1C0 \sr_60_[2]  (.D(\sr_59_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_60_[2]_net_1 ));
    DFN1E1C0 \sr_26_[7]  (.D(\sr_25_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_26_[7]_net_1 ));
    DFN1E1C0 \sr_2_[0]  (.D(sr_prev[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_5), .Q(\sr_2_[0]_net_1 ));
    DFN1E1C0 \sr_41_[9]  (.D(\sr_40_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_41_[9]_net_1 ));
    DFN1E1C0 \sr_57_[0]  (.D(\sr_56_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_57_[0]_net_1 ));
    DFN1E1C0 \sr_48_[8]  (.D(\sr_47_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_48_[8]_net_1 ));
    DFN1E1C0 \sr_53_[1]  (.D(\sr_52_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_53_[1]_net_1 ));
    DFN1E1C0 \sr_2_[6]  (.D(sr_prev[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_5), .Q(\sr_2_[6]_net_1 ));
    DFN1E1C0 \sr_7_[7]  (.D(\sr_6_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_7_[7]_net_1 ));
    DFN1E1C0 \sr_42_[1]  (.D(\sr_41_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_42_[1]_net_1 ));
    DFN1E1C0 \sr_63_[1]  (.D(\sr_62_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[1]));
    DFN1E1C0 \sr_50_[4]  (.D(\sr_49_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_50_[4]_net_1 ));
    DFN1E1C0 \sr_58_[12]  (.D(\sr_57_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_58_[12]_net_1 ));
    DFN1E1C0 \sr_58_[3]  (.D(\sr_57_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_58_[3]_net_1 ));
    DFN1E1C0 \sr_28_[2]  (.D(\sr_27_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_28_[2]_net_1 ));
    DFN1E1C0 \sr_4_[2]  (.D(\sr_3_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_4_[2]_net_1 ));
    DFN1E1C0 \sr_4_[8]  (.D(\sr_3_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_4_[8]_net_1 ));
    DFN1E1C0 \sr_28_[5]  (.D(\sr_27_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_28_[5]_net_1 ));
    DFN1E1C0 \sr_28_[12]  (.D(\sr_27_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_28_[12]_net_1 ));
    DFN1E1C0 \sr_60_[4]  (.D(\sr_59_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_60_[4]_net_1 ));
    DFN1E1C0 \sr_19_[11]  (.D(\sr_18_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_19_[11]_net_1 ));
    DFN1E1C0 \sr_14_[9]  (.D(\sr_13_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_14_[9]_net_1 ));
    DFN1E1C0 \sr_18_[8]  (.D(\sr_17_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_18_[8]_net_1 ));
    DFN1E1C0 \sr_47_[11]  (.D(\sr_46_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_47_[11]_net_1 ));
    DFN1E1C0 \sr_20_[7]  (.D(\sr_19_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_20_[7]_net_1 ));
    DFN1E1C0 \sr_2_[1]  (.D(sr_prev[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_5), .Q(\sr_2_[1]_net_1 ));
    DFN1E1C0 \sr_31_[0]  (.D(\sr_30_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_31_[0]_net_1 ));
    DFN1E1C0 \sr_42_[10]  (.D(\sr_41_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_42_[10]_net_1 ));
    DFN1E1C0 \sr_44_[0]  (.D(\sr_43_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_44_[0]_net_1 ));
    DFN1E1C0 \sr_13_[7]  (.D(\sr_12_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_13_[7]_net_1 ));
    DFN1E1C0 \sr_36_[12]  (.D(\sr_35_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_36_[12]_net_1 ));
    DFN1E1C0 \sr_9_[5]  (.D(\sr_8_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[5]_net_1 ));
    DFN1E1C0 \sr_34_[12]  (.D(\sr_33_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_34_[12]_net_1 ));
    DFN1E1C0 \sr_3_[7]  (.D(\sr_2_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_3_[7]_net_1 ));
    DFN1E1C0 \sr_13_[6]  (.D(\sr_12_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_13_[6]_net_1 ));
    DFN1E1C0 \sr_16_[9]  (.D(\sr_15_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_16_[9]_net_1 ));
    DFN1E1C0 \sr_12_[12]  (.D(\sr_11_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_12_[12]_net_1 ));
    DFN1E1C0 \sr_43_[5]  (.D(\sr_42_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_43_[5]_net_1 ));
    DFN1E1C0 \sr_46_[0]  (.D(\sr_45_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_46_[0]_net_1 ));
    DFN1E1C0 \sr_52_[2]  (.D(\sr_51_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_52_[2]_net_1 ));
    DFN1E1C0 \sr_60_[9]  (.D(\sr_59_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_60_[9]_net_1 ));
    DFN1E1C0 \sr_4_[12]  (.D(\sr_3_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_4_[12]_net_1 ));
    DFN1E1C0 \sr_58_[11]  (.D(\sr_57_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_58_[11]_net_1 ));
    DFN1E1C0 \sr_3_[12]  (.D(\sr_2_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_3_[12]_net_1 ));
    DFN1E1C0 \sr_23_[9]  (.D(\sr_22_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_23_[9]_net_1 ));
    DFN1E1C0 \sr_28_[11]  (.D(\sr_27_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_28_[11]_net_1 ));
    DFN1E1C0 \sr_62_[2]  (.D(\sr_61_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_62_[2]_net_1 ));
    DFN1E1C0 \sr_16_[11]  (.D(\sr_15_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_16_[11]_net_1 ));
    DFN1E1C0 \sr_1_[12]  (.D(sr_new_0_0), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_27), .Q(sr_prev[12]));
    DFN1E1C0 \sr_18_[2]  (.D(\sr_17_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_18_[2]_net_1 ));
    DFN1E1C0 \sr_39_[1]  (.D(\sr_38_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_39_[1]_net_1 ));
    DFN1E1C0 \sr_23_[1]  (.D(\sr_22_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_23_[1]_net_1 ));
    DFN1E1C0 \sr_18_[0]  (.D(\sr_17_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_18_[0]_net_1 ));
    DFN1E1C0 \sr_38_[8]  (.D(\sr_37_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[8]_net_1 ));
    DFN1E1C0 \sr_8_[10]  (.D(\sr_7_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_8_[10]_net_1 ));
    DFN1E1C0 \sr_10_[9]  (.D(\sr_9_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_10_[9]_net_1 ));
    DFN1E1C0 \sr_45_[12]  (.D(\sr_44_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_45_[12]_net_1 ));
    DFN1E1C0 \sr_39_[2]  (.D(\sr_38_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_39_[2]_net_1 ));
    DFN1E1C0 \sr_8_[12]  (.D(\sr_7_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_8_[12]_net_1 ));
    DFN1E1C0 \sr_15_[11]  (.D(\sr_14_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_15_[11]_net_1 ));
    DFN1E1C0 \sr_39_[7]  (.D(\sr_38_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_39_[7]_net_1 ));
    DFN1E1C0 \sr_52_[4]  (.D(\sr_51_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_52_[4]_net_1 ));
    DFN1E1C0 \sr_41_[4]  (.D(\sr_40_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_41_[4]_net_1 ));
    DFN1E1C0 \sr_58_[5]  (.D(\sr_57_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_58_[5]_net_1 ));
    DFN1E1C0 \sr_40_[0]  (.D(\sr_39_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_40_[0]_net_1 ));
    DFN1E1C0 \sr_31_[3]  (.D(\sr_30_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_31_[3]_net_1 ));
    DFN1E1C0 \sr_51_[6]  (.D(\sr_50_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_51_[6]_net_1 ));
    DFN1E1C0 \sr_17_[12]  (.D(\sr_16_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_17_[12]_net_1 ));
    DFN1E1C0 \sr_45_[3]  (.D(\sr_44_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_45_[3]_net_1 ));
    DFN1E1C0 \sr_62_[4]  (.D(\sr_61_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_62_[4]_net_1 ));
    DFN1E1C0 \sr_21_[4]  (.D(\sr_20_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_21_[4]_net_1 ));
    DFN1E1C0 \sr_60_[3]  (.D(\sr_59_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_60_[3]_net_1 ));
    DFN1E1C0 \sr_22_[7]  (.D(\sr_21_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_22_[7]_net_1 ));
    DFN1E1C0 \sr_61_[6]  (.D(\sr_60_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_61_[6]_net_1 ));
    DFN1E1C0 \sr_49_[9]  (.D(\sr_48_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_49_[9]_net_1 ));
    DFN1E1C0 \sr_18_[10]  (.D(\sr_17_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_18_[10]_net_1 ));
    DFN1E1C0 \sr_8_[5]  (.D(\sr_7_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_8_[5]_net_1 ));
    DFN1E1C0 \sr_33_[12]  (.D(\sr_32_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_33_[12]_net_1 ));
    DFN1E1C0 \sr_28_[3]  (.D(\sr_27_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_28_[3]_net_1 ));
    DFN1E1C0 \sr_38_[9]  (.D(\sr_37_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[9]_net_1 ));
    DFN1E1C0 \sr_53_[11]  (.D(\sr_52_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_53_[11]_net_1 ));
    DFN1E1C0 \sr_37_[1]  (.D(\sr_36_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[1]_net_1 ));
    DFN1E1C0 \sr_37_[2]  (.D(\sr_36_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[2]_net_1 ));
    DFN1E1C0 \sr_23_[11]  (.D(\sr_22_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_23_[11]_net_1 ));
    DFN1E1C0 \sr_3_[11]  (.D(\sr_2_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_3_[11]_net_1 ));
    DFN1E1C0 \sr_37_[7]  (.D(\sr_36_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[7]_net_1 ));
    DFN1E1C0 \sr_38_[6]  (.D(\sr_37_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[6]_net_1 ));
    DFN1E1C0 \sr_41_[6]  (.D(\sr_40_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_41_[6]_net_1 ));
    DFN1E1C0 \sr_44_[7]  (.D(\sr_43_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_44_[7]_net_1 ));
    DFN1E1C0 \sr_54_[7]  (.D(\sr_53_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_54_[7]_net_1 ));
    DFN1E1C0 \sr_0_[7]  (.D(cur_error[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_21), .Q(sr_new[7]));
    DFN1E1C0 \sr_9_[11]  (.D(\sr_8_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_9_[11]_net_1 ));
    DFN1E1C0 \sr_62_[9]  (.D(\sr_61_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_62_[9]_net_1 ));
    DFN1E1C0 \sr_54_[8]  (.D(\sr_53_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_54_[8]_net_1 ));
    DFN1E1C0 \sr_39_[0]  (.D(\sr_38_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_39_[0]_net_1 ));
    DFN1E1C0 \sr_47_[9]  (.D(\sr_46_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_47_[9]_net_1 ));
    DFN1E1C0 \sr_6_[12]  (.D(\sr_5_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_6_[12]_net_1 ));
    DFN1E1C0 \sr_7_[11]  (.D(\sr_6_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_7_[11]_net_1 ));
    DFN1E1C0 \sr_46_[7]  (.D(\sr_45_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_46_[7]_net_1 ));
    DFN1E1C0 \sr_14_[5]  (.D(\sr_13_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_14_[5]_net_1 ));
    DFN1E1C0 \sr_56_[7]  (.D(\sr_55_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_56_[7]_net_1 ));
    DFN1E1C0 \sr_12_[9]  (.D(\sr_11_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_12_[9]_net_1 ));
    DFN1E1C0 \sr_12_[11]  (.D(\sr_11_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_12_[11]_net_1 ));
    DFN1E1C0 \sr_55_[9]  (.D(\sr_54_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_55_[9]_net_1 ));
    DFN1E1C0 \sr_56_[8]  (.D(\sr_55_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_56_[8]_net_1 ));
    DFN1E1C0 \sr_25_[6]  (.D(\sr_24_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_25_[6]_net_1 ));
    DFN1E1C0 \sr_14_[3]  (.D(\sr_13_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_14_[3]_net_1 ));
    DFN1E1C0 \sr_42_[0]  (.D(\sr_41_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_42_[0]_net_1 ));
    DFN1E1C0 \sr_1_[7]  (.D(sr_new[7]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable_31), .Q(sr_prev[7]));
    DFN1E1C0 \sr_2_[5]  (.D(sr_prev[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_5), .Q(\sr_2_[5]_net_1 ));
    DFN1E1C0 \sr_14_[11]  (.D(\sr_13_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_14_[11]_net_1 ));
    DFN1E1C0 \sr_37_[0]  (.D(\sr_36_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_37_[0]_net_1 ));
    DFN1E1C0 \sr_58_[1]  (.D(\sr_57_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_58_[1]_net_1 ));
    DFN1E1C0 \sr_11_[1]  (.D(\sr_10_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_11_[1]_net_1 ));
    DFN1E1C0 \sr_62_[3]  (.D(\sr_61_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_62_[3]_net_1 ));
    DFN1E1C0 \sr_45_[10]  (.D(\sr_44_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_45_[10]_net_1 ));
    DFN1E1C0 \sr_16_[5]  (.D(\sr_15_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_16_[5]_net_1 ));
    DFN1E1C0 \sr_43_[3]  (.D(\sr_42_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_43_[3]_net_1 ));
    DFN1E1C0 \sr_61_[5]  (.D(\sr_60_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_61_[5]_net_1 ));
    DFN1E1C0 \sr_54_[0]  (.D(\sr_53_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_54_[0]_net_1 ));
    DFN1E1C0 \sr_16_[3]  (.D(\sr_15_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_16_[3]_net_1 ));
    DFN1E1C0 \sr_4_[9]  (.D(\sr_3_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_4_[9]_net_1 ));
    DFN1E1C0 \sr_40_[7]  (.D(\sr_39_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_40_[7]_net_1 ));
    DFN1E1C0 \sr_50_[7]  (.D(\sr_49_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_50_[7]_net_1 ));
    DFN1E1C0 \sr_31_[5]  (.D(\sr_30_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_31_[5]_net_1 ));
    DFN1E1C0 \sr_50_[8]  (.D(\sr_49_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_50_[8]_net_1 ));
    DFN1E1C0 \sr_49_[4]  (.D(\sr_48_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_49_[4]_net_1 ));
    DFN1E1C0 \sr_31_[4]  (.D(\sr_30_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_31_[4]_net_1 ));
    DFN1E1C0 \sr_0_[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable_5), .Q(sr_new[12]));
    DFN1E1C0 \sr_39_[3]  (.D(\sr_38_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_39_[3]_net_1 ));
    DFN1E1C0 \sr_6_[7]  (.D(\sr_5_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_6_[7]_net_1 ));
    DFN1E1C0 \sr_60_[7]  (.D(\sr_59_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_60_[7]_net_1 ));
    DFN1E1C0 \sr_59_[6]  (.D(\sr_58_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_59_[6]_net_1 ));
    DFN1E1C0 \sr_7_[3]  (.D(\sr_6_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_7_[3]_net_1 ));
    DFN1E1C0 \sr_46_[10]  (.D(\sr_45_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_46_[10]_net_1 ));
    DFN1E1C0 \sr_60_[8]  (.D(\sr_59_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_60_[8]_net_1 ));
    DFN1E1C0 \sr_29_[4]  (.D(\sr_28_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(\sr_29_[4]_net_1 ));
    DFN1E1C0 \sr_57_[11]  (.D(\sr_56_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_5), .Q(\sr_57_[11]_net_1 ));
    DFN1E1C0 \sr_56_[0]  (.D(\sr_55_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_56_[0]_net_1 ));
    DFN1E1C0 \sr_5_[7]  (.D(\sr_4_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_5_[7]_net_1 ));
    DFN1E1C0 \sr_18_[7]  (.D(\sr_17_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_18_[7]_net_1 ));
    DFN1E1C0 \sr_10_[5]  (.D(\sr_9_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_10_[5]_net_1 ));
    DFN1E1C0 \sr_41_[12]  (.D(\sr_40_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_41_[12]_net_1 ));
    DFN1E1C0 \sr_52_[10]  (.D(\sr_51_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_52_[10]_net_1 ));
    DFN1E1C0 \sr_27_[11]  (.D(\sr_26_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_27_[11]_net_1 ));
    DFN1E1C0 \sr_39_[12]  (.D(\sr_38_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_39_[12]_net_1 ));
    DFN1E1C0 \sr_18_[6]  (.D(\sr_17_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_18_[6]_net_1 ));
    DFN1E1C0 \sr_22_[10]  (.D(\sr_21_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_22_[10]_net_1 ));
    DFN1E1C0 \sr_10_[3]  (.D(\sr_9_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_10_[3]_net_1 ));
    DFN1E1C0 \sr_48_[5]  (.D(\sr_47_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_48_[5]_net_1 ));
    DFN1E1C0 \sr_60_[0]  (.D(\sr_59_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_60_[0]_net_1 ));
    DFN1E1C0 \sr_47_[4]  (.D(\sr_46_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_47_[4]_net_1 ));
    DFN1E1C0 \sr_30_[12]  (.D(\sr_29_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_30_[12]_net_1 ));
    DFN1E1C0 \sr_37_[3]  (.D(\sr_36_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[3]_net_1 ));
    DFN1E1C0 \sr_57_[6]  (.D(\sr_56_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_57_[6]_net_1 ));
    DFN1E1C0 \sr_49_[6]  (.D(\sr_48_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_49_[6]_net_1 ));
    DFN1E1C0 \sr_3_[3]  (.D(\sr_2_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_3_[3]_net_1 ));
    DFN1E1C0 \sr_28_[9]  (.D(\sr_27_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_28_[9]_net_1 ));
    DFN1E1C0 \sr_27_[4]  (.D(\sr_26_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_27_[4]_net_1 ));
    DFN1E1C0 \sr_62_[12]  (.D(\sr_61_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_62_[12]_net_1 ));
    DFN1E1C0 \sr_50_[0]  (.D(\sr_49_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_50_[0]_net_1 ));
    DFN1E1C0 \sr_53_[9]  (.D(\sr_52_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_53_[9]_net_1 ));
    DFN1E1C0 \sr_23_[6]  (.D(\sr_22_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_23_[6]_net_1 ));
    DFN1E1C0 \sr_28_[1]  (.D(\sr_27_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_28_[1]_net_1 ));
    DFN1E1C0 \sr_11_[4]  (.D(\sr_10_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_11_[4]_net_1 ));
    DFN1E1C0 \sr_30_[10]  (.D(\sr_29_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_30_[10]_net_1 ));
    DFN1E1C0 \sr_21_[8]  (.D(\sr_20_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_21_[8]_net_1 ));
    DFN1E1C0 \sr_16_[12]  (.D(\sr_15_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_16_[12]_net_1 ));
    DFN1E1C0 \sr_41_[10]  (.D(\sr_40_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_41_[10]_net_1 ));
    DFN1E1C0 \sr_45_[1]  (.D(\sr_44_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_45_[1]_net_1 ));
    DFN1E1C0 \sr_33_[10]  (.D(\sr_32_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_33_[10]_net_1 ));
    DFN1E1C0 \sr_14_[12]  (.D(\sr_13_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_14_[12]_net_1 ));
    DFN1E1C0 \sr_41_[11]  (.D(\sr_40_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_41_[11]_net_1 ));
    DFN1E1C0 \sr_55_[12]  (.D(\sr_54_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_55_[12]_net_1 ));
    DFN1E1C0 \sr_42_[7]  (.D(\sr_41_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_42_[7]_net_1 ));
    DFN1E1C0 \sr_52_[7]  (.D(\sr_51_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_52_[7]_net_1 ));
    DFN1E1C0 \sr_41_[2]  (.D(\sr_40_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_41_[2]_net_1 ));
    DFN1E1C0 \sr_52_[8]  (.D(\sr_51_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_52_[8]_net_1 ));
    DFN1E1C0 \sr_25_[12]  (.D(\sr_24_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_25_[12]_net_1 ));
    DFN1E1C0 \sr_47_[6]  (.D(\sr_46_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_47_[6]_net_1 ));
    DFN1E1C0 \sr_62_[7]  (.D(\sr_61_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_62_[7]_net_1 ));
    DFN1E1C0 \sr_62_[8]  (.D(\sr_61_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_62_[8]_net_1 ));
    DFN1E1C0 \sr_19_[1]  (.D(\sr_18_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_19_[1]_net_1 ));
    DFN1E1C0 \sr_21_[0]  (.D(\sr_20_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_21_[0]_net_1 ));
    DFN1E1C0 \sr_39_[10]  (.D(\sr_38_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_39_[10]_net_1 ));
    DFN1E1C0 \sr_12_[5]  (.D(\sr_11_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_12_[5]_net_1 ));
    DFN1E1C0 \sr_0_[10]  (.D(cur_error[10]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable_5), .Q(sr_new[10]));
    DFN1E1C0 \sr_12_[3]  (.D(\sr_11_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_12_[3]_net_1 ));
    DFN1E1C0 \sr_34_[1]  (.D(\sr_33_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_34_[1]_net_1 ));
    DFN1E1C0 \sr_39_[5]  (.D(\sr_38_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_39_[5]_net_1 ));
    DFN1E1C0 \sr_5_[11]  (.D(\sr_4_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_5_[11]_net_1 ));
    DFN1E1C0 \sr_34_[2]  (.D(\sr_33_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_34_[2]_net_1 ));
    DFN1E1C0 \sr_39_[4]  (.D(\sr_38_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_39_[4]_net_1 ));
    DFN1E1C0 \sr_55_[2]  (.D(\sr_54_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_55_[2]_net_1 ));
    DFN1E1C0 \sr_62_[0]  (.D(\sr_61_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_62_[0]_net_1 ));
    DFN1E1C0 \sr_34_[7]  (.D(\sr_33_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_34_[7]_net_1 ));
    DFN1E1C0 \sr_41_[8]  (.D(\sr_40_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_41_[8]_net_1 ));
    DFN1E1C0 \sr_52_[0]  (.D(\sr_51_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_52_[0]_net_1 ));
    DFN1E1C0 \sr_17_[1]  (.D(\sr_16_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_17_[1]_net_1 ));
    DFN1E1C0 \sr_4_[0]  (.D(\sr_3_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_4_[0]_net_1 ));
    DFN1E1C0 \sr_36_[1]  (.D(\sr_35_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_36_[1]_net_1 ));
    DFN1E1C0 \sr_13_[12]  (.D(\sr_12_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_13_[12]_net_1 ));
    DFN1E1C0 \sr_4_[6]  (.D(\sr_3_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_4_[6]_net_1 ));
    DFN1E1C0 \sr_44_[9]  (.D(\sr_43_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_44_[9]_net_1 ));
    DFN1E1C0 \sr_0_[3]  (.D(cur_error[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_21), .Q(sr_new[3]));
    DFN1E1C0 \sr_36_[2]  (.D(\sr_35_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_36_[2]_net_1 ));
    DFN1E1C0 \sr_51_[3]  (.D(\sr_50_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_51_[3]_net_1 ));
    DFN1E1C0 \sr_36_[7]  (.D(\sr_35_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_36_[7]_net_1 ));
    DFN1E1C0 \sr_21_[2]  (.D(\sr_20_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_21_[2]_net_1 ));
    DFN1E1C0 \sr_37_[5]  (.D(\sr_36_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[5]_net_1 ));
    DFN1E1C0 \sr_55_[4]  (.D(\sr_54_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_55_[4]_net_1 ));
    DFN1E1C0 \sr_21_[5]  (.D(\sr_20_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_21_[5]_net_1 ));
    DFN1E1C0 \sr_43_[1]  (.D(\sr_42_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_43_[1]_net_1 ));
    DFN1E1C0 \sr_11_[8]  (.D(\sr_10_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_11_[8]_net_1 ));
    DFN1E1C0 \sr_37_[4]  (.D(\sr_36_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[4]_net_1 ));
    DFN1E1C0 \sr_62_[11]  (.D(\sr_61_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_62_[11]_net_1 ));
    DFN1E1C0 \sr_46_[9]  (.D(\sr_45_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_46_[9]_net_1 ));
    DFN1E1C0 \sr_25_[7]  (.D(\sr_24_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_25_[7]_net_1 ));
    DFN1E1C0 \sr_48_[3]  (.D(\sr_47_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_48_[3]_net_1 ));
    DFN1E1C0 \sr_30_[1]  (.D(\sr_29_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_30_[1]_net_1 ));
    DFN1E1C0 \sr_4_[1]  (.D(\sr_3_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_4_[1]_net_1 ));
    DFN1E1C0 \sr_55_[10]  (.D(\sr_54_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(\sr_55_[10]_net_1 ));
    DFN1E1C0 \sr_19_[4]  (.D(\sr_18_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_19_[4]_net_1 ));
    DFN1E1C0 \sr_9_[7]  (.D(\sr_8_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[7]_net_1 ));
    DFN1E1C0 \sr_7_[4]  (.D(\sr_6_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_7_[4]_net_1 ));
    DFN1E1C0 \sr_29_[8]  (.D(\sr_28_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(\sr_29_[8]_net_1 ));
    DFN1E1C0 \sr_1_[3]  (.D(sr_new[3]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable_30), .Q(sr_prev[3]));
    DFN1E1C0 \sr_34_[0]  (.D(\sr_33_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_34_[0]_net_1 ));
    DFN1E1C0 \sr_30_[2]  (.D(\sr_29_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_30_[2]_net_1 ));
    DFN1E1C0 \sr_25_[10]  (.D(\sr_24_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_25_[10]_net_1 ));
    DFN1E1C0 \sr_30_[7]  (.D(\sr_29_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_30_[7]_net_1 ));
    DFN1E1C0 \sr_49_[2]  (.D(\sr_48_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_49_[2]_net_1 ));
    DFN1E1C0 \sr_56_[10]  (.D(\sr_55_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_56_[10]_net_1 ));
    DFN1E1C0 \sr_40_[9]  (.D(\sr_39_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_40_[9]_net_1 ));
    DFN1E1C0 \sr_36_[0]  (.D(\sr_35_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_36_[0]_net_1 ));
    DFN1E1C0 \sr_11_[2]  (.D(\sr_10_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_11_[2]_net_1 ));
    DFN1E1C0 \sr_30_[11]  (.D(\sr_29_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_30_[11]_net_1 ));
    DFN1E1C0 \sr_53_[2]  (.D(\sr_52_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_53_[2]_net_1 ));
    DFN1E1C0 \sr_26_[10]  (.D(\sr_25_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_26_[10]_net_1 ));
    DFN1E1C0 \sr_11_[0]  (.D(\sr_10_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_11_[0]_net_1 ));
    DFN1E1C0 \sr_31_[8]  (.D(\sr_30_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_31_[8]_net_1 ));
    DFN1E1C0 \sr_29_[0]  (.D(\sr_28_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_29_[0]_net_1 ));
    DFN1E1C0 \sr_17_[4]  (.D(\sr_16_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_17_[4]_net_1 ));
    DFN1E1C0 \sr_6_[3]  (.D(\sr_5_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_6_[3]_net_1 ));
    DFN1E1C0 \sr_51_[12]  (.D(\sr_50_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_51_[12]_net_1 ));
    DFN1E1C0 \sr_27_[8]  (.D(\sr_26_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_27_[8]_net_1 ));
    DFN1E1C0 \sr_3_[4]  (.D(\sr_2_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_3_[4]_net_1 ));
    DFN1E1C0 \sr_63_[2]  (.D(\sr_62_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[2]));
    DFN1E1C0 \sr_21_[12]  (.D(\sr_20_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_21_[12]_net_1 ));
    DFN1E1C0 \sr_5_[3]  (.D(\sr_4_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_5_[3]_net_1 ));
    DFN1E1C0 \sr_15_[9]  (.D(\sr_14_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_15_[9]_net_1 ));
    DFN1E1C0 \sr_51_[5]  (.D(\sr_50_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_51_[5]_net_1 ));
    DFN1E1C0 \sr_47_[2]  (.D(\sr_46_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_47_[2]_net_1 ));
    DFN1E1C0 \sr_47_[10]  (.D(\sr_46_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_47_[10]_net_1 ));
    DFN1E1C0 \sr_45_[0]  (.D(\sr_44_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_45_[0]_net_1 ));
    DFN1E1C0 \sr_58_[9]  (.D(\sr_57_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_58_[9]_net_1 ));
    DFN1E1C0 \sr_30_[0]  (.D(\sr_29_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_30_[0]_net_1 ));
    DFN1E1C0 \sr_44_[4]  (.D(\sr_43_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_44_[4]_net_1 ));
    DFN1E1C0 \sr_53_[4]  (.D(\sr_52_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_53_[4]_net_1 ));
    DFN1E1C0 \sr_34_[3]  (.D(\sr_33_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_34_[3]_net_1 ));
    DFN1E1C0 \sr_54_[6]  (.D(\sr_53_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_54_[6]_net_1 ));
    DFN1E1C0 \sr_49_[8]  (.D(\sr_48_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_49_[8]_net_1 ));
    DFN1E1C0 \sr_28_[6]  (.D(\sr_27_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_19), .Q(\sr_28_[6]_net_1 ));
    DFN1E1C0 \sr_21_[3]  (.D(\sr_20_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_21_[3]_net_1 ));
    DFN1E1C0 \sr_31_[9]  (.D(\sr_30_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_31_[9]_net_1 ));
    DFN1E1C0 \sr_8_[7]  (.D(\sr_7_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_8_[7]_net_1 ));
    DFN1E1C0 \sr_27_[0]  (.D(\sr_26_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_27_[0]_net_1 ));
    DFN1E1C0 \sr_24_[4]  (.D(\sr_23_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_24_[4]_net_1 ));
    DFN1E1C0 \sr_63_[4]  (.D(\sr_62_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[4]));
    DFN1E1C0 \sr_32_[1]  (.D(\sr_31_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_32_[1]_net_1 ));
    DFN1E1C0 \sr_19_[12]  (.D(\sr_18_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_19_[12]_net_1 ));
    DFN1E1C0 \sr_23_[7]  (.D(\sr_22_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_23_[7]_net_1 ));
    DFN1E1C0 \sr_51_[10]  (.D(\sr_50_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_51_[10]_net_1 ));
    DFN1E1C0 \sr_32_[2]  (.D(\sr_31_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_32_[2]_net_1 ));
    DFN1E1C0 \sr_38_[12]  (.D(\sr_37_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[12]_net_1 ));
    DFN1E1C0 \sr_59_[3]  (.D(\sr_58_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_59_[3]_net_1 ));
    DFN1E1C0 \sr_51_[11]  (.D(\sr_50_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_51_[11]_net_1 ));
    DFN1E1C0 \sr_29_[2]  (.D(\sr_28_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(\sr_29_[2]_net_1 ));
    DFN1E1C0 \sr_32_[7]  (.D(\sr_31_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_32_[7]_net_1 ));
    DFN1E1C0 \sr_21_[10]  (.D(\sr_20_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_21_[10]_net_1 ));
    DFN1E1C0 \sr_46_[4]  (.D(\sr_45_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_46_[4]_net_1 ));
    DFN1E1C0 \sr_31_[6]  (.D(\sr_30_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_31_[6]_net_1 ));
    DFN1E1C0 \sr_36_[3]  (.D(\sr_35_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_24), .Q(\sr_36_[3]_net_1 ));
    DFN1E1C0 \sr_29_[5]  (.D(\sr_28_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(\sr_29_[5]_net_1 ));
    DFN1E1C0 \sr_56_[6]  (.D(\sr_55_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_56_[6]_net_1 ));
    DFN1E1C0 \sr_21_[11]  (.D(\sr_20_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_21_[11]_net_1 ));
    DFN1E1C0 \sr_19_[8]  (.D(\sr_18_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_19_[8]_net_1 ));
    DFN1E1C0 \sr_44_[10]  (.D(\sr_43_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_32), .Q(\sr_44_[10]_net_1 ));
    DFN1E1C0 \sr_10_[12]  (.D(\sr_9_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_10_[12]_net_1 ));
    DFN1E1C0 \sr_26_[4]  (.D(\sr_25_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_26_[4]_net_1 ));
    DFN1E1C0 \sr_47_[8]  (.D(\sr_46_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_20), .Q(\sr_47_[8]_net_1 ));
    DFN1E1C0 \sr_44_[6]  (.D(\sr_43_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_28), .Q(\sr_44_[6]_net_1 ));
    DFN1E1C0 \sr_42_[9]  (.D(\sr_41_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_42_[9]_net_1 ));
    DFN1E1C0 \sr_63_[9]  (.D(\sr_62_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[9]));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \sr_10_[10]  (.D(\sr_9_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_10_[10]_net_1 ));
    DFN1E1C0 \sr_2_[10]  (.D(sr_prev[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_14), .Q(\sr_2_[10]_net_1 ));
    DFN1E1C0 \sr_13_[10]  (.D(\sr_12_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_13_[10]_net_1 ));
    DFN1E1C0 \sr_57_[3]  (.D(\sr_56_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_9), .Q(\sr_57_[3]_net_1 ));
    DFN1E1C0 \sr_27_[2]  (.D(\sr_26_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_27_[2]_net_1 ));
    DFN1E1C0 \sr_40_[4]  (.D(\sr_39_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_40_[4]_net_1 ));
    DFN1E1C0 \sr_30_[3]  (.D(\sr_29_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_30_[3]_net_1 ));
    DFN1E1C0 \sr_50_[6]  (.D(\sr_49_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_50_[6]_net_1 ));
    DFN1E1C0 \sr_27_[5]  (.D(\sr_26_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_27_[5]_net_1 ));
    DFN1E1C0 \sr_46_[6]  (.D(\sr_45_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_12), .Q(\sr_46_[6]_net_1 ));
    DFN1E1C0 \sr_38_[11]  (.D(\sr_37_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_38_[11]_net_1 ));
    DFN1E1C0 \sr_17_[8]  (.D(\sr_16_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_17_[8]_net_1 ));
    DFN1E1C0 \sr_20_[4]  (.D(\sr_19_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_20_[4]_net_1 ));
    DFN1E1C0 \sr_0_[4]  (.D(cur_error[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_21), .Q(sr_new[4]));
    DFN1E1C0 \sr_49_[11]  (.D(\sr_48_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_49_[11]_net_1 ));
    DFN1E1C0 \sr_13_[9]  (.D(\sr_12_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_21), .Q(\sr_13_[9]_net_1 ));
    DFN1E1C0 \sr_60_[6]  (.D(\sr_59_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_2), .Q(\sr_60_[6]_net_1 ));
    DFN1E1C0 \sr_2_[7]  (.D(sr_prev[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable_5), .Q(\sr_2_[7]_net_1 ));
    DFN1E1C0 \sr_51_[1]  (.D(\sr_50_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_51_[1]_net_1 ));
    DFN1E1C0 \sr_32_[0]  (.D(\sr_31_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_32_[0]_net_1 ));
    DFN1E1C0 \sr_7_[2]  (.D(\sr_6_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_15), .Q(\sr_7_[2]_net_1 ));
    DFN1E1C0 \sr_4_[11]  (.D(\sr_3_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_4_[11]_net_1 ));
    DFN1E1C0 \sr_19_[2]  (.D(\sr_18_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_19_[2]_net_1 ));
    DFN1E1C0 \sr_7_[8]  (.D(\sr_6_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_16), .Q(\sr_7_[8]_net_1 ));
    DFN1E1C0 \sr_4_[5]  (.D(\sr_3_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_4_[5]_net_1 ));
    DFN1E1C0 \sr_43_[0]  (.D(\sr_42_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_18), .Q(\sr_43_[0]_net_1 ));
    DFN1E1C0 \sr_19_[0]  (.D(\sr_18_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_7), .Q(\sr_19_[0]_net_1 ));
    DFN1E1C0 \sr_9_[10]  (.D(\sr_8_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_33), .Q(\sr_9_[10]_net_1 ));
    DFN1E1C0 \sr_39_[8]  (.D(\sr_38_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_39_[8]_net_1 ));
    DFN1E1C0 \sr_61_[1]  (.D(\sr_60_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_11), .Q(\sr_61_[1]_net_1 ));
    DFN1E1C0 \sr_19_[10]  (.D(\sr_18_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_10), .Q(\sr_19_[10]_net_1 ));
    DFN1E1C0 \sr_14_[1]  (.D(\sr_13_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_31), .Q(\sr_14_[1]_net_1 ));
    DFN1E1C0 \sr_63_[3]  (.D(\sr_62_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[3]));
    DFN1E1C0 \sr_45_[7]  (.D(\sr_44_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_3), .Q(\sr_45_[7]_net_1 ));
    DFN1E1C0 \sr_59_[5]  (.D(\sr_58_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_27), .Q(\sr_59_[5]_net_1 ));
    DFN1E1C0 \sr_55_[7]  (.D(\sr_54_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_55_[7]_net_1 ));
    DFN1E1C0 \sr_63_[12]  (.D(\sr_62_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(sr_old[12]));
    DFN1E1C0 \sr_48_[1]  (.D(\sr_47_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_30), .Q(\sr_48_[1]_net_1 ));
    DFN1E1C0 \sr_42_[12]  (.D(\sr_41_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_22), .Q(\sr_42_[12]_net_1 ));
    DFN1E1C0 \sr_40_[6]  (.D(\sr_39_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_26), .Q(\sr_40_[6]_net_1 ));
    DFN1E1C0 \sr_55_[8]  (.D(\sr_54_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_25), .Q(\sr_55_[8]_net_1 ));
    DFN1E1C0 \sr_1_[4]  (.D(sr_new[4]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable_30), .Q(sr_prev[4]));
    DFN1E1C0 \sr_34_[5]  (.D(\sr_33_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_34_[5]_net_1 ));
    DFN1E1C0 \sr_6_[11]  (.D(\sr_5_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_1), .Q(\sr_6_[11]_net_1 ));
    DFN1E1C0 \sr_11_[7]  (.D(\sr_10_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_11_[7]_net_1 ));
    DFN1E1C0 \sr_34_[4]  (.D(\sr_33_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_6), .Q(\sr_34_[4]_net_1 ));
    DFN1E1C0 \sr_16_[1]  (.D(\sr_15_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_14), .Q(\sr_16_[1]_net_1 ));
    DFN1E1C0 \sr_29_[3]  (.D(\sr_28_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_29), .Q(\sr_29_[3]_net_1 ));
    DFN1E1C0 \sr_17_[2]  (.D(\sr_16_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_17_[2]_net_1 ));
    DFN1E1C0 \sr_39_[9]  (.D(\sr_38_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_17), .Q(\sr_39_[9]_net_1 ));
    DFN1E1C0 \sr_3_[2]  (.D(\sr_2_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_3_[2]_net_1 ));
    DFN1E1C0 \sr_46_[11]  (.D(\sr_45_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_8), .Q(\sr_46_[11]_net_1 ));
    DFN1E1C0 \sr_3_[8]  (.D(\sr_2_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_13), .Q(\sr_3_[8]_net_1 ));
    DFN1E1C0 \sr_33_[11]  (.D(\sr_32_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_0), .Q(\sr_33_[11]_net_1 ));
    DFN1E1C0 \sr_17_[0]  (.D(\sr_16_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_23), .Q(\sr_17_[0]_net_1 ));
    DFN1E1C0 \sr_37_[8]  (.D(\sr_36_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[8]_net_1 ));
    DFN1E1C0 \sr_15_[5]  (.D(\sr_14_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_5), .Q(\sr_15_[5]_net_1 ));
    DFN1E1C0 \sr_11_[6]  (.D(\sr_10_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable_4), .Q(\sr_11_[6]_net_1 ));
    
endmodule


module controller_Z1_4_1(
       state_0_d0,
       state_0_0,
       pwm_chg,
       int_done,
       sig_prev,
       sig_old_i_0,
       avg_done,
       int_enable,
       vd_rdy,
       sum_rdy,
       deriv_enable,
       calc_avg,
       calc_int,
       pwm_enable,
       sum_enable,
       avg_enable,
       pwm_chg_0,
       int_enable_0,
       int_enable_1,
       int_enable_2,
       int_enable_3,
       int_enable_4,
       int_enable_5,
       int_enable_6,
       int_enable_7,
       int_enable_8,
       int_enable_9,
       int_enable_10,
       int_enable_11,
       int_enable_12,
       int_enable_13,
       int_enable_14,
       int_enable_15,
       int_enable_16,
       int_enable_17,
       int_enable_18,
       int_enable_19,
       int_enable_20,
       int_enable_21,
       int_enable_22,
       int_enable_23,
       int_enable_24,
       int_enable_25,
       int_enable_26,
       int_enable_27,
       int_enable_28,
       int_enable_29,
       int_enable_30,
       int_enable_31,
       int_enable_32,
       int_enable_33,
       avg_enable_0,
       n_rst_c,
       clk_c,
       avg_enable_1,
       calc_error
    );
input  state_0_d0;
input  state_0_0;
output pwm_chg;
input  int_done;
input  sig_prev;
input  sig_old_i_0;
input  avg_done;
output int_enable;
input  vd_rdy;
input  sum_rdy;
output deriv_enable;
output calc_avg;
output calc_int;
output pwm_enable;
output sum_enable;
output avg_enable;
output pwm_chg_0;
output int_enable_0;
output int_enable_1;
output int_enable_2;
output int_enable_3;
output int_enable_4;
output int_enable_5;
output int_enable_6;
output int_enable_7;
output int_enable_8;
output int_enable_9;
output int_enable_10;
output int_enable_11;
output int_enable_12;
output int_enable_13;
output int_enable_14;
output int_enable_15;
output int_enable_16;
output int_enable_17;
output int_enable_18;
output int_enable_19;
output int_enable_20;
output int_enable_21;
output int_enable_22;
output int_enable_23;
output int_enable_24;
output int_enable_25;
output int_enable_26;
output int_enable_27;
output int_enable_28;
output int_enable_29;
output int_enable_30;
output int_enable_31;
output int_enable_32;
output int_enable_33;
output avg_enable_0;
input  n_rst_c;
input  clk_c;
output avg_enable_1;
output calc_error;

    wire N_170_0, \state[7]_net_1 , N_24, \state_RNI6K7H2[0]_net_1 , 
        \state_RNIHDCF1_0[7]_net_1 , N_12, N_94, count_31_0, count_c13, 
        count_n14, \count[14]_net_1 , N_62, count_n13, count_c12, 
        \count[13]_net_1 , count_n11, count_c10, \count[11]_net_1 , 
        count_n12, count_c11, \count[12]_net_1 , count_n15, 
        \count[15]_net_1 , count_c7, count_c6, \count[7]_net_1 , 
        count_c5, \count[6]_net_1 , count_c4, \count[5]_net_1 , 
        count_c3, \count[4]_net_1 , count_c2, \count[3]_net_1 , 
        count_c1, \count[2]_net_1 , \count[0]_net_1 , \count[1]_net_1 , 
        count_c8, \count[8]_net_1 , count_c9, \count[9]_net_1 , 
        \count[10]_net_1 , \state_ns_0_a2_9[0] , \state[10]_net_1 , 
        N_33, \state_ns_0_a2_8[0] , \state_ns_0_a2_6[0] , 
        \state_ns_0_a2_5[0] , \state_ns_0_a2_2[0] , N_270, 
        \state_RNIH6UI_0[12]_net_1 , \state_ns_0_a2_1[0] , 
        \state_ns_0_a2_0[0] , next_state_0_sqmuxa_1_1_a2_0_a2_0, 
        \state_ns_i_0_0[2] , un1_countlto15_13, un1_countlto15_5, 
        un1_countlto15_4, un1_countlto15_11, un1_countlto15_12, 
        un1_countlto15_1, un1_countlto15_0, un1_countlto15_9, 
        un1_countlto15_7, un1_countlto15_3, N_274, N_273, 
        \state[0]_net_1 , N_26, next_state15_li, 
        \state_RNI4V7Q[4]_net_1 , N_23, count_n7, count_n6, count_n5, 
        count_n4, count_n3, count_n2, count_n8, count_n9, count_n10, 
        \state[4]_net_1 , \state[12]_net_1 , \avg_count[0]_net_1 , 
        \avg_count[1]_net_1 , N_27, \state_ns[1] , \state_ns[0] , 
        \state_ns[12] , \state_ns[10] , \state_ns[4] , count_n1, N_267, 
        counte, \state_RNO_1[8] , \state_ns[7] , 
        \DWACT_ADD_CI_0_partial_sum[0] , I_10_1, 
        \DWACT_ADD_CI_0_TMP[0] , GND, VCC;
    
    DFN1C0 \state_11[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_11));
    DFN1P0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .PRE(n_rst_c), 
        .Q(\state[0]_net_1 ));
    DFN1E1C0 \count[15]  (.D(count_n15), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[15]_net_1 ));
    XA1B \count_RNO[6]  (.A(\count[6]_net_1 ), .B(count_c5), .C(N_62), 
        .Y(count_n6));
    XA1B \count_RNO[3]  (.A(\count[3]_net_1 ), .B(count_c2), .C(N_62), 
        .Y(count_n3));
    NOR2B \count_RNI4ABH3[7]  (.A(count_c6), .B(\count[7]_net_1 ), .Y(
        count_c7));
    DFN1E1C0 \count[9]  (.D(count_n9), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[9]_net_1 ));
    AO1A \state_RNO[10]  (.A(sum_rdy), .B(\state[10]_net_1 ), .C(
        sum_enable), .Y(\state_ns[10] ));
    OR2A \state_RNIC8TE[7]  (.A(vd_rdy), .B(\state[7]_net_1 ), .Y(
        \state_ns_i_0_0[2] ));
    DFN1C0 \state_1[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_1));
    NOR2 \state_RNO_6[0]  (.A(sum_enable), .B(\state[7]_net_1 ), .Y(
        \state_ns_0_a2_2[0] ));
    DFN1C0 \state[10]  (.D(\state_ns[10] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[10]_net_1 ));
    DFN1C0 \state_0[13]  (.D(N_12), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_chg_0));
    DFN1E1C0 \count[8]  (.D(count_n8), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[8]_net_1 ));
    XA1B \count_RNO[1]  (.A(\count[1]_net_1 ), .B(\count[0]_net_1 ), 
        .C(N_62), .Y(count_n1));
    DFN1C0 \state_21[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_21));
    DFN1C0 \state[6]  (.D(int_enable), .CLK(clk_c), .CLR(n_rst_c), .Q(
        calc_int));
    XA1B \count_RNO[12]  (.A(count_c11), .B(\count[12]_net_1 ), .C(
        N_62), .Y(count_n12));
    DFN1C0 \state_4[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_4));
    DFN1C0 \state_0[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_0));
    OR2 \state_RNO[12]  (.A(N_27), .B(pwm_enable), .Y(\state_ns[12] ));
    XA1B \count_RNO[2]  (.A(\count[2]_net_1 ), .B(count_c1), .C(N_62), 
        .Y(count_n2));
    XA1B \count_RNO[11]  (.A(count_c10), .B(\count[11]_net_1 ), .C(
        N_62), .Y(count_n11));
    AND2 un1_avg_count_1_I_1 (.A(\avg_count[0]_net_1 ), .B(
        \state_RNI4V7Q[4]_net_1 ), .Y(\DWACT_ADD_CI_0_TMP[0] ));
    DFN1E1C0 \count[10]  (.D(count_n10), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[10]_net_1 ));
    DFN1C0 \state_32[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_32));
    DFN1E1C0 \count[5]  (.D(count_n5), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[5]_net_1 ));
    NOR2 \count_RNIDMAS[1]  (.A(\count[2]_net_1 ), .B(\count[1]_net_1 )
        , .Y(un1_countlto15_1));
    DFN1C0 \state[4]  (.D(\state_ns[4] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[4]_net_1 ));
    NOR2B \state_RNI4V7Q[4]  (.A(\state[4]_net_1 ), .B(avg_done), .Y(
        \state_RNI4V7Q[4]_net_1 ));
    NOR2B \count_RNI20GA1[2]  (.A(count_c1), .B(\count[2]_net_1 ), .Y(
        count_c2));
    DFN1C0 \state_30[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_30));
    DFN1C0 \state[7]  (.D(\state_ns[7] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[7]_net_1 ));
    AO1 \state_RNIISGR5[10]  (.A(sig_old_i_0), .B(sig_prev), .C(N_62), 
        .Y(counte));
    DFN1C0 \state[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable));
    DFN1E1C0 \count[4]  (.D(count_n4), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[4]_net_1 ));
    GND GND_i (.Y(GND));
    NOR3A \state_RNIS6S51[0]  (.A(N_273), .B(\state[10]_net_1 ), .C(
        \state[0]_net_1 ), .Y(N_274));
    DFN1C0 \state_15[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_15));
    DFN1E1C0 \count[12]  (.D(count_n12), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[12]_net_1 ));
    DFN1E1C0 \count[0]  (.D(N_267), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[0]_net_1 ));
    DFN1C0 \avg_count[1]  (.D(I_10_1), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \avg_count[1]_net_1 ));
    DFN1C0 \state_12[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_12));
    XA1B \count_RNO[5]  (.A(\count[5]_net_1 ), .B(count_c4), .C(N_62), 
        .Y(count_n5));
    NOR2 \count_RNILUAS[5]  (.A(\count[6]_net_1 ), .B(\count[5]_net_1 )
        , .Y(un1_countlto15_3));
    XOR2 un1_avg_count_1_I_8 (.A(\avg_count[0]_net_1 ), .B(
        \state_RNI4V7Q[4]_net_1 ), .Y(\DWACT_ADD_CI_0_partial_sum[0] ));
    NOR2 \count_RNIJHT6[13]  (.A(\count[14]_net_1 ), .B(
        \count[13]_net_1 ), .Y(un1_countlto15_7));
    AX1 \count_RNO[15]  (.A(N_62), .B(\count[15]_net_1 ), .C(N_94), .Y(
        count_n15));
    NOR2B \count_RNIVEMD4[9]  (.A(count_c8), .B(\count[9]_net_1 ), .Y(
        count_c9));
    NOR2A \state_RNO[1]  (.A(\state_RNI4V7Q[4]_net_1 ), .B(
        next_state15_li), .Y(\state_ns[1] ));
    DFN1C0 \state_19[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_19));
    DFN1C0 \state_10[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_10));
    DFN1C0 \state_25[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_25));
    OA1A \state_RNO_0[0]  (.A(\state[10]_net_1 ), .B(N_33), .C(
        \state_ns_0_a2_8[0] ), .Y(\state_ns_0_a2_9[0] ));
    DFN1C0 \state_18[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_18));
    DFN1C0 \state_22[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_22));
    NOR2A \state_RNIF8CS[10]  (.A(\state_RNIH6UI_0[12]_net_1 ), .B(
        \state[10]_net_1 ), .Y(N_24));
    DFN1C0 \state[12]  (.D(\state_ns[12] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[12]_net_1 ));
    VCC VCC_i (.Y(VCC));
    NOR3A \state_RNIHDCF1_0[7]  (.A(calc_error), .B(\state[7]_net_1 ), 
        .C(N_24), .Y(\state_RNIHDCF1_0[7]_net_1 ));
    NOR2 \state_RNIU4ES[0]  (.A(\state_RNIH6UI_0[12]_net_1 ), .B(
        \state[0]_net_1 ), .Y(N_23));
    XA1B \count_RNO[14]  (.A(count_c13), .B(\count[14]_net_1 ), .C(
        N_62), .Y(count_n14));
    DFN1E1C0 \count[13]  (.D(count_n13), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[13]_net_1 ));
    AO1A \state_RNO[4]  (.A(avg_done), .B(\state[4]_net_1 ), .C(
        calc_avg), .Y(\state_ns[4] ));
    DFN1C0 \state_29[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_29));
    DFN1C0 \state_20[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_20));
    XOR2 un1_avg_count_1_I_10 (.A(\avg_count[1]_net_1 ), .B(
        \DWACT_ADD_CI_0_TMP[0] ), .Y(I_10_1));
    DFN1C0 \state[9]  (.D(deriv_enable), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(sum_enable));
    OR2B \avg_count_RNI5AKA[1]  (.A(\avg_count[0]_net_1 ), .B(
        \avg_count[1]_net_1 ), .Y(next_state15_li));
    NOR2 \count_RNI48KH[10]  (.A(\count[9]_net_1 ), .B(
        \count[10]_net_1 ), .Y(un1_countlto15_5));
    DFN1C0 \state_28[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_28));
    NOR2 \count_RNO[0]  (.A(\count[0]_net_1 ), .B(N_62), .Y(N_267));
    NOR2 \count_RNIP2BS[7]  (.A(\count[7]_net_1 ), .B(\count[8]_net_1 )
        , .Y(un1_countlto15_4));
    NOR3B \state_RNO_3[0]  (.A(\state_ns_0_a2_6[0] ), .B(
        \state_ns_0_a2_5[0] ), .C(avg_enable), .Y(\state_ns_0_a2_8[0] )
        );
    DFN1C0 \state_16[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_16));
    DFN1E1C0 \count[1]  (.D(count_n1), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[1]_net_1 ));
    XA1B \count_RNO[7]  (.A(\count[7]_net_1 ), .B(count_c6), .C(N_62), 
        .Y(count_n7));
    DFN1E1C0 \count[3]  (.D(count_n3), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[3]_net_1 ));
    NOR2B \count_RNO_0[15]  (.A(count_31_0), .B(count_c13), .Y(N_94));
    XA1B \count_RNO[9]  (.A(count_c8), .B(\count[9]_net_1 ), .C(N_62), 
        .Y(count_n9));
    AO1A \state_RNO[7]  (.A(int_done), .B(\state[7]_net_1 ), .C(
        calc_int), .Y(\state_ns[7] ));
    AOI1B \state_RNIEVII5[10]  (.A(un1_countlto15_13), .B(
        un1_countlto15_12), .C(next_state_0_sqmuxa_1_1_a2_0_a2_0), .Y(
        N_62));
    DFN1C0 \state[13]  (.D(N_12), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_chg));
    NOR3A \count_RNI2VQD[11]  (.A(un1_countlto15_7), .B(
        \count[12]_net_1 ), .C(\count[11]_net_1 ), .Y(
        un1_countlto15_11));
    DFN1C0 \state_7[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_7));
    DFN1C0 \avg_count[0]  (.D(\DWACT_ADD_CI_0_partial_sum[0] ), .CLK(
        clk_c), .CLR(n_rst_c), .Q(\avg_count[0]_net_1 ));
    DFN1C0 \state[8]  (.D(\state_RNO_1[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(deriv_enable));
    DFN1C0 \state_26[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_26));
    DFN1C0 \state_14[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_14));
    NOR2B \count_RNICQJK4[11]  (.A(count_c10), .B(\count[11]_net_1 ), 
        .Y(count_c11));
    OR2B \state_RNIH6UI[12]  (.A(\state[4]_net_1 ), .B(
        \state[12]_net_1 ), .Y(N_273));
    DFN1C0 \state[3]  (.D(avg_enable), .CLK(clk_c), .CLR(n_rst_c), .Q(
        calc_avg));
    NOR3C \count_RNIJJK63[15]  (.A(un1_countlto15_1), .B(
        un1_countlto15_0), .C(un1_countlto15_9), .Y(un1_countlto15_12));
    XA1B \count_RNO[4]  (.A(\count[4]_net_1 ), .B(count_c3), .C(N_62), 
        .Y(count_n4));
    XA1B \count_RNO[13]  (.A(count_c12), .B(\count[13]_net_1 ), .C(
        N_62), .Y(count_n13));
    DFN1C0 \state_2[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_2));
    NOR2B \count_RNIQCLO1[3]  (.A(count_c2), .B(\count[3]_net_1 ), .Y(
        count_c3));
    NOR3A \count_RNI6PLO1[3]  (.A(un1_countlto15_3), .B(
        \count[3]_net_1 ), .C(\count[4]_net_1 ), .Y(un1_countlto15_9));
    NOR2B \count_RNI8P533[6]  (.A(count_c5), .B(\count[6]_net_1 ), .Y(
        count_c6));
    NOR3B \state_RNO_5[0]  (.A(\state_ns_0_a2_1[0] ), .B(
        \state_ns_0_a2_0[0] ), .C(calc_error), .Y(\state_ns_0_a2_5[0] )
        );
    NOR2B \count_RNIKH2O4[12]  (.A(count_c11), .B(\count[12]_net_1 ), 
        .Y(count_c12));
    DFN1C0 \state_24[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_24));
    DFN1C0 \state_8[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_8));
    DFN1C0 \state_1[2]  (.D(\state_RNI6K7H2[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable_1));
    NOR2 \state_RNO_8[0]  (.A(pwm_enable), .B(calc_int), .Y(
        \state_ns_0_a2_1[0] ));
    NOR3B \state_RNO_1[0]  (.A(next_state15_li), .B(
        \state_RNI4V7Q[4]_net_1 ), .C(\state[10]_net_1 ), .Y(N_26));
    NOR3B \state_RNO_4[0]  (.A(\state_ns_0_a2_2[0] ), .B(N_270), .C(
        \state_RNIH6UI_0[12]_net_1 ), .Y(\state_ns_0_a2_6[0] ));
    NOR2B \count_RNIBKAS[1]  (.A(\count[0]_net_1 ), .B(
        \count[1]_net_1 ), .Y(count_c1));
    NOR3C \count_RNIV9QR1[10]  (.A(un1_countlto15_5), .B(
        un1_countlto15_4), .C(un1_countlto15_11), .Y(un1_countlto15_13)
        );
    NOR2 \count_RNI04KH[15]  (.A(\count[15]_net_1 ), .B(
        \count[0]_net_1 ), .Y(un1_countlto15_0));
    DFN1E1C0 \count[7]  (.D(count_n7), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[7]_net_1 ));
    DFN1C0 \state[2]  (.D(\state_RNI6K7H2[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable));
    DFN1C0 \state_33[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_33));
    DFN1C0 \state_0[2]  (.D(\state_RNI6K7H2[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable_0));
    DFN1C0 \state_6[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_6));
    DFN1C0 \state_17[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_17));
    DFN1C0 \state[1]  (.D(\state_ns[1] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(calc_error));
    DFN1E1C0 \count[6]  (.D(count_n6), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[6]_net_1 ));
    OA1 \state_RNO_0[12]  (.A(state_0_0), .B(state_0_d0), .C(
        \state[12]_net_1 ), .Y(N_27));
    NOR2B \count_RNI1SGV3[8]  (.A(count_c7), .B(\count[8]_net_1 ), .Y(
        count_c8));
    DFN1C0 \state_5[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_5));
    DFN1C0 \state_3[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_3));
    NOR2B \state_RNO[8]  (.A(\state[7]_net_1 ), .B(int_done), .Y(
        \state_RNO_1[8] ));
    AO1A \state_RNO[0]  (.A(int_enable), .B(\state_ns_0_a2_9[0] ), .C(
        N_26), .Y(\state_ns[0] ));
    NOR2B \count_RNIT9HR4[13]  (.A(count_c12), .B(\count[13]_net_1 ), 
        .Y(count_c13));
    DFN1C0 \state_9[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_9));
    NOR2B \count_RNID90L2[5]  (.A(count_c4), .B(\count[5]_net_1 ), .Y(
        count_c5));
    OR2 \state_RNIH6UI_0[12]  (.A(\state[4]_net_1 ), .B(
        \state[12]_net_1 ), .Y(\state_RNIH6UI_0[12]_net_1 ));
    NOR3C \state_RNO_2[0]  (.A(un1_countlto15_12), .B(
        un1_countlto15_13), .C(sum_rdy), .Y(N_33));
    NOR3A \state_RNIHDCF1[7]  (.A(calc_error), .B(\state[7]_net_1 ), 
        .C(N_24), .Y(N_170_0));
    DFN1C0 \state_27[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_27));
    DFN1C0 \state[11]  (.D(N_62), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_enable));
    DFN1E1C0 \count[2]  (.D(count_n2), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[2]_net_1 ));
    NOR3A \state_RNIV0011[12]  (.A(\state[12]_net_1 ), .B(state_0_0), 
        .C(state_0_d0), .Y(N_12));
    DFN1C0 \state_31[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_31));
    NOR2 \state_RNO_9[0]  (.A(calc_avg), .B(deriv_enable), .Y(
        \state_ns_0_a2_0[0] ));
    XA1B \count_RNO[8]  (.A(count_c7), .B(\count[8]_net_1 ), .C(N_62), 
        .Y(count_n8));
    NOR2B \state_RNIS14G[10]  (.A(\state[10]_net_1 ), .B(sum_rdy), .Y(
        next_state_0_sqmuxa_1_1_a2_0_a2_0));
    DFN1C0 \state_13[5]  (.D(\state_RNIHDCF1_0[7]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(int_enable_13));
    NOR2B \count_RNI545H4[10]  (.A(count_c9), .B(\count[10]_net_1 ), 
        .Y(count_c10));
    DFN1E1C0 \count[11]  (.D(count_n11), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[11]_net_1 ));
    NOR3 \state_RNI6K7H2[0]  (.A(N_274), .B(\state_ns_i_0_0[2] ), .C(
        N_23), .Y(\state_RNI6K7H2[0]_net_1 ));
    NOR2A \count_RNO_1[15]  (.A(\count[14]_net_1 ), .B(N_62), .Y(
        count_31_0));
    NOR2B \count_RNIJQQ62[4]  (.A(count_c3), .B(\count[4]_net_1 ), .Y(
        count_c4));
    DFN1E1C0 \count[14]  (.D(count_n14), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[14]_net_1 ));
    XA1B \count_RNO[10]  (.A(count_c9), .B(\count[10]_net_1 ), .C(N_62)
        , .Y(count_n10));
    OR2B \state_RNO_7[0]  (.A(vd_rdy), .B(\state[0]_net_1 ), .Y(N_270));
    DFN1C0 \state_23[5]  (.D(N_170_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        int_enable_23));
    
endmodule


module sig_gen_4(
       primary_fb_c,
       n_rst_c,
       clk_c,
       sig_old_i_0,
       sig_prev
    );
input  primary_fb_c;
input  n_rst_c;
input  clk_c;
output sig_old_i_0;
output sig_prev;

    wire sig_prev_i, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(clk_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev_inst_1 (.D(primary_fb_c), .CLK(clk_c), .CLR(
        n_rst_c), .Q(sig_prev));
    INV sig_old_RNO (.A(sig_prev), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module pid_sum_13s_4_1(
       integral_i,
       integral,
       sr_new,
       derivative_0,
       sr_new_1_0,
       sr_new_0_0,
       integral_1_0,
       integral_0_0,
       sum_39,
       sum_14,
       sum_20,
       sum_19,
       sum_22,
       sum_13,
       sum_17,
       sum_18,
       sum_21,
       sum_23,
       sum_16,
       sum_15,
       sum_12,
       sum_11,
       sum_6,
       sum_10,
       sum_9,
       sum_5,
       sum_8,
       sum_7,
       sum_4,
       sum_2_d0,
       sum_1_d0,
       sum_0_d0,
       sum_3,
       sum_0_0,
       sum_1_0,
       sum_2_0,
       sum_enable,
       sum_rdy,
       n_rst_c,
       clk_c
    );
input  [25:24] integral_i;
input  [25:6] integral;
input  [12:0] sr_new;
input  derivative_0;
input  sr_new_1_0;
input  sr_new_0_0;
input  integral_1_0;
input  integral_0_0;
output sum_39;
output sum_14;
output sum_20;
output sum_19;
output sum_22;
output sum_13;
output sum_17;
output sum_18;
output sum_21;
output sum_23;
output sum_16;
output sum_15;
output sum_12;
output sum_11;
output sum_6;
output sum_10;
output sum_9;
output sum_5;
output sum_8;
output sum_7;
output sum_4;
output sum_2_d0;
output sum_1_d0;
output sum_0_d0;
output sum_3;
output sum_0_0;
output sum_1_0;
output sum_2_0;
input  sum_enable;
output sum_rdy;
input  n_rst_c;
input  clk_c;

    wire \next_sum[39] , \state_RNI172K[6]_net_1 , \state_0[1]_net_1 , 
        \state_RNIK76G[0]_net_1 , \state_2[2]_net_1 , 
        \state_1[2]_net_1 , \state_0[2]_net_1 , \state_0[3]_net_1 , 
        \state[6]_net_1 , N_416_0, \un1_next_sum_1_iv_0[26] , 
        next_sum_1_sqmuxa_2, next_sum_1_sqmuxa_1, next_sum_1_sqmuxa, 
        N_12, N_10, \DWACT_FINC_E[0] , N_5, \DWACT_FINC_E[4] , N_2, 
        \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , N_25, N_23, 
        \DWACT_FINC_E_0[0] , N_18, \DWACT_FINC_E_0[4] , N_15, 
        \DWACT_FINC_E_0[7] , \DWACT_FINC_E_0[6] , 
        ADD_40x40_fast_I448_Y_0, \sumreg[30]_net_1 , 
        \un1_next_sum_1_iv[26] , ADD_40x40_fast_I447_Y_0, 
        \sumreg[29]_net_1 , ADD_40x40_fast_I456_Y_0, 
        \sumreg[38]_net_1 , ADD_40x40_fast_I449_Y_0, 
        \sumreg[31]_net_1 , ADD_40x40_fast_I453_Y_0, 
        \sumreg[35]_net_1 , ADD_40x40_fast_I454_Y_0, 
        \sumreg[36]_net_1 , ADD_40x40_fast_I455_Y_0, 
        \sumreg[37]_net_1 , ADD_40x40_fast_I452_Y_0, 
        \sumreg[34]_net_1 , ADD_40x40_fast_I451_Y_0, 
        \sumreg[33]_net_1 , ADD_40x40_fast_I347_Y_0, N787, N772, N771, 
        ADD_40x40_fast_I457_Y_0, ADD_40x40_fast_I446_Y_0, 
        \sumreg[28]_net_1 , ADD_40x40_fast_I450_Y_0, 
        \sumreg[32]_net_1 , ADD_40x40_fast_I348_Y_0, N789, N774, N773, 
        ADD_40x40_fast_I379_Y_3, N756, ADD_40x40_fast_I379_Y_2, N596, 
        ADD_40x40_fast_I379_Y_0, N681, ADD_40x40_fast_I346_Y_0, N785, 
        N770, N769, ADD_40x40_fast_I382_Y_2, I274_un1_Y, 
        ADD_40x40_fast_I382_Y_0, I382_un1_Y, N679, N687, 
        ADD_40x40_fast_I381_Y_2, N760, N775, ADD_40x40_fast_I381_Y_1, 
        N600, N685, ADD_40x40_fast_I445_Y_0, \sumreg[27]_net_1 , 
        ADD_40x40_fast_I380_Y_3, I270_un1_Y, ADD_40x40_fast_I380_Y_1, 
        I380_un1_Y, I122_un1_Y, N594, N683, ADD_40x40_fast_I432_Y_0, 
        \un1_next_sum_iv_1[14] , \un1_next_sum_iv_2[14] , 
        ADD_40x40_fast_I438_Y_0, \un1_next_sum[20] , 
        ADD_40x40_fast_I437_Y_0, \un1_next_sum[19] , 
        ADD_40x40_fast_I347_un1_Y_0, N788, ADD_40x40_fast_I384_Y_2, 
        ADD_40x40_fast_I384_un1_Y_0, N850, ADD_40x40_fast_I384_Y_1, 
        N766, N781, ADD_40x40_fast_I384_Y_0, N691, N684, 
        ADD_40x40_fast_I383_Y_2, ADD_40x40_fast_I383_un1_Y_0, N848, 
        ADD_40x40_fast_I383_Y_1, N764, N779, ADD_40x40_fast_I383_Y_0, 
        N689, ADD_40x40_fast_I444_Y_0, \sumreg[26]_net_1 , 
        ADD_40x40_fast_I443_Y_0, \sumreg[25]_net_1 , 
        \un1_next_sum_0_iv[25] , ADD_40x40_fast_I440_Y_0, 
        \un1_next_sum[22] , ADD_40x40_fast_I378_Y_3, N754, 
        ADD_40x40_fast_I378_Y_2, ADD_40x40_fast_I378_Y_0, 
        ADD_40x40_fast_I431_Y_0, \un1_next_sum_iv_1[13] , 
        \un1_next_sum_iv_2[13] , ADD_40x40_fast_I349_Y_0, N791, N776, 
        ADD_40x40_fast_I435_Y_0, \un1_next_sum_iv_1[17] , 
        \un1_next_sum_iv_2[17] , ADD_40x40_fast_I436_Y_0, 
        \un1_next_sum_iv_1[18] , \un1_next_sum_iv_2[18] , 
        ADD_40x40_fast_I385_Y_2, I280_un1_Y, ADD_40x40_fast_I385_Y_0, 
        I385_un1_Y, N693, N686, ADD_40x40_fast_I442_Y_0, 
        \sumreg[24]_net_1 , \un1_next_sum[24] , 
        ADD_40x40_fast_I348_un1_Y_0, N790, ADD_40x40_fast_I439_Y_0, 
        \un1_next_sum[21] , ADD_40x40_fast_I441_Y_0, 
        \un1_next_sum[23] , ADD_40x40_fast_I434_Y_0, 
        \un1_next_sum_iv_1[16] , \un1_next_sum_iv_2[16] , 
        ADD_40x40_fast_I433_Y_0, \un1_next_sum_iv_1[15] , 
        \un1_next_sum_iv_2[15] , ADD_40x40_fast_I346_un1_Y_0, N786, 
        ADD_40x40_fast_I350_Y_0, N793, N778, N777, 
        ADD_40x40_fast_I351_Y_0, I292_un1_Y, ADD_40x40_fast_I430_Y_0, 
        \un1_next_sum_iv_1[12] , \un1_next_sum_iv_2[12] , 
        ADD_40x40_fast_I349_un1_Y_0, N792, ADD_40x40_fast_I353_Y_0, 
        N799, N784, N783, ADD_40x40_fast_I429_Y_0, 
        \un1_next_sum_iv_1[11] , \un1_next_sum_iv_2[11] , 
        ADD_40x40_fast_I350_un1_Y_0, N794, ADD_40x40_fast_I424_Y_0, 
        \un1_next_sum[6] , ADD_40x40_fast_I428_Y_0, 
        \un1_next_sum_iv_1[10] , \un1_next_sum_iv_2[10] , 
        ADD_40x40_fast_I427_Y_0, \un1_next_sum[9] , 
        ADD_40x40_fast_I351_un1_Y_0, N706, N698, N796, 
        ADD_40x40_fast_I352_un1_Y_0, N798, N782, 
        ADD_40x40_fast_I423_Y_0, \un1_next_sum[5] , 
        ADD_40x40_fast_I426_Y_0, \un1_next_sum_iv_1[8] , 
        \un1_next_sum_iv_2[8] , ADD_40x40_fast_I353_un1_Y_0, N800, 
        ADD_40x40_fast_I425_Y_0, \un1_next_sum_iv_1[7] , 
        \un1_next_sum_iv_2[7] , N814, N666, N812, N745, 
        ADD_40x40_fast_I422_Y_0, \un1_next_sum[4] , 
        ADD_40x40_fast_I420_Y_0, \un1_next_sum[0] , 
        ADD_40x40_fast_I419_Y_0, ADD_40x40_fast_I257_Y_1, N475, N472, 
        N661, ADD_40x40_fast_I195_Y_0, ADD_40x40_fast_I197_Y_0, 
        ADD_40x40_fast_I187_Y_0, ADD_22x22_fast_I126_Y_1, N371, N378, 
        ADD_22x22_fast_I126_Y_0, N335, N332, N331, 
        ADD_22x22_fast_I142_Y_0_1, ADD_22x22_fast_I142_Y_0_a3_0, N329, 
        ADD_22x22_fast_I142_Y_0_0, \i_adj[18]_net_1 , 
        \i_adj[20]_net_1 , N_14_1, ADD_22x22_fast_I172_Y_0, 
        \i_adj[12]_net_1 , \i_adj[14]_net_1 , 
        ADD_22x22_fast_I126_un1_Y_0, N379, 
        ADD_22x22_fast_I142_Y_0_a3_1, N330, ADD_40x40_fast_I418_Y_0, 
        ADD_22x22_fast_I177_Y_0, \i_adj[19]_net_1 , \i_adj[17]_net_1 , 
        ADD_22x22_fast_I178_Y_0, ADD_40x40_fast_I421_Y_0, N743, 
        ADD_22x22_fast_I130_Y_0, N386, ADD_22x22_fast_I142_Y_0_o3_0_0, 
        N337, N334, N333, ADD_22x22_fast_I143_Y_3, 
        ADD_22x22_fast_I143_un1_Y_0, N423, ADD_22x22_fast_I143_Y_2, 
        N367, N374, ADD_22x22_fast_I143_Y_1, N328, 
        ADD_22x22_fast_I143_Y_0, N314, ADD_22x22_fast_I144_Y_2, 
        ADD_22x22_fast_I144_un1_Y_0, N425, ADD_22x22_fast_I144_Y_1, 
        N369, N376, ADD_22x22_fast_I144_Y_0, \un1_next_sum_iv_0[20] , 
        \ireg[20]_net_1 , \un1_next_sum_iv_0[21] , \ireg[21]_net_1 , 
        \un1_next_sum_iv_0[23] , \ireg[23]_net_1 , 
        \un1_next_sum_iv_0[4] , \ireg[4]_net_1 , 
        \un1_next_sum_iv_0[5] , \ireg[5]_net_1 , 
        \un1_next_sum_iv_0[22] , \ireg[22]_net_1 , 
        \un1_next_sum_iv_0[19] , \ireg[19]_net_1 , 
        \un1_next_sum_iv_0[24] , \ireg[24]_net_1 , 
        ADD_22x22_fast_I128_Y_0, N382, N375, ADD_22x22_fast_I170_Y_0, 
        \i_adj[10]_net_1 , ADD_22x22_fast_I169_Y_0, \i_adj[9]_net_1 , 
        \i_adj[11]_net_1 , \un24_next_sum_m[16] , next_sum_0_sqmuxa_1, 
        \un3_next_sum_m[16] , \preg[16]_net_1 , \ireg_m[16] , 
        \un24_next_sum_m[8] , \un3_next_sum_m[8] , \preg[8]_net_1 , 
        \ireg_m[8] , \un1_next_sum_iv_2[6] , \un24_next_sum_m[6] , 
        \un3_next_sum_m[6] , \un1_next_sum_iv_1[6] , \preg[6]_net_1 , 
        \ireg_m[6] , \un24_next_sum_m[7] , \un3_next_sum_m[7] , 
        \preg[7]_net_1 , \ireg_m[7] , \un24_next_sum_m[13] , 
        \un3_next_sum_m[13] , \preg[13]_net_1 , \ireg_m[13] , 
        \un24_next_sum_m[12] , \un3_next_sum_m[12] , \preg[12]_net_1 , 
        \ireg_m[12] , \un24_next_sum_m[15] , \un3_next_sum_m[15] , 
        \preg[15]_net_1 , \ireg_m[15] , \un1_next_sum_iv_2[9] , 
        \un24_next_sum_m[9] , \un3_next_sum_m[9] , 
        \un1_next_sum_iv_1[9] , \preg[9]_net_1 , \ireg_m[9] , 
        \un24_next_sum_m[17] , \un3_next_sum_m[17] , \preg[17]_net_1 , 
        \ireg_m[17] , \un24_next_sum_m[10] , \un3_next_sum_m[10] , 
        \preg[10]_net_1 , \ireg_m[10] , \un24_next_sum_m[11] , 
        \un3_next_sum_m[11] , \preg[11]_net_1 , \ireg_m[11] , 
        \un24_next_sum_m[14] , \un3_next_sum_m[14] , \preg[14]_net_1 , 
        \ireg_m[14] , \un24_next_sum_m[18] , \un3_next_sum_m[18] , 
        \preg[18]_net_1 , \ireg_m[18] , ADD_22x22_fast_I142_Y_0_a3_3_0, 
        N338, ADD_m8_i_1, next_sum_0_sqmuxa_2, ADD_m8_i_a4_0_1, 
        \un1_next_sum_0_iv_1[25] , \un3_next_sum_m[25] , 
        ADD_22x22_fast_I129_Y_0, N384, N377, ADD_22x22_fast_I166_Y_0, 
        \i_adj[6]_net_1 , \i_adj[8]_net_1 , 
        ADD_22x22_fast_I128_un1_Y_0, N383, ADD_22x22_fast_I131_Y_0, 
        N345, N342, N341, ADD_22x22_fast_I165_Y_0, \i_adj[7]_net_1 , 
        \i_adj[5]_net_1 , ADD_22x22_fast_I129_un1_Y_0, N385, N266, 
        N359, ADD_22x22_fast_I163_Y_0, \i_adj[3]_net_1 , N_9, 
        ADD_22x22_fast_I85_Y_0, \i_adj[2]_net_1 , \i_adj[4]_net_1 , 
        N270, ADD_m8_i_a4_0_0, ADD_m8_i_o4_1, ADD_m8_i_a4_4, N_232, 
        N492, N_11, N393, N354, \next_ireg_3[15] , N424, I133_un1_Y, 
        \next_ireg_3[7] , \i_adj[1]_net_1 , \next_ireg_3[9] , N396, 
        \next_ireg_3[25] , \i_adj[21]_net_1 , N1049, N1097, N1031, 
        N879, \next_ireg_3[11] , N531, N1029, N846, N877, N878, N1027, 
        I381_un1_Y, I336_un1_Y, N876, N823, N844, N597, N601, N884, 
        N852, N1035, N883, N1040, N1088, N595, N680, I378_un1_Y, N817, 
        N870, N838, N1021, I330_un1_Y, N1033, N881, \next_ireg_3[23] , 
        I124_un1_Y, \next_ireg_3[8] , \next_ireg_3[10] , N394, 
        \next_ireg_3[16] , N422, I132_un1_Y, \next_ireg_3[13] , N525, 
        \next_ireg_3[19] , \i_adj[13]_net_1 , \i_adj[15]_net_1 , N507, 
        \next_ireg_3[20] , \i_adj[16]_net_1 , N504, \next_ireg_3[21] , 
        \next_ireg_3[22] , N498, \next_ireg_3[24] , I122_un1_Y_0, 
        \next_ireg_3[18] , I130_un1_Y, \next_ireg_3[17] , N513, 
        \next_ireg_3[14] , N522, \next_ireg_3[12] , N528, 
        \state[5]_net_1 , \state[4]_net_1 , next_sum_0_sqmuxa, 
        \ireg_m[25] , N1025, N842, N873, N821, N874, N1023, I332_un1_Y, 
        I379_un1_Y, N840, N872, N819, N1058, N1106, N1055, I294_un1_Y, 
        I352_un1_Y, N1103, N1052, N1100, N1046, N1094, N1043, N1091, 
        N1037, N1085, N758, N599, N682, N816, N734, I131_un1_Y, 
        I106_un1_Y, N389, N381, N387, \state[1]_net_1 , N740, N659, 
        \inf_abs1_5[0] , \inf_abs1_5[3] , \inf_abs1_a_2[3] , 
        \inf_abs1_5[12] , \inf_abs1_a_2[12] , \inf_abs1_5[1] , 
        \inf_abs1_a_2[1] , \inf_abs1_5[2] , \inf_abs1_a_2[2] , 
        \inf_abs1_5[4] , \inf_abs1_a_2[4] , \inf_abs1_5[6] , 
        \inf_abs1_a_2[6] , \inf_abs1_5[9] , \inf_abs1_a_2[9] , 
        \inf_abs1_5[11] , \inf_abs1_a_2[11] , \state[3]_net_1 , 
        \ireg[17]_net_1 , \next_sum[18] , N1076, I359_un1_Y, 
        \inf_abs2_5[3] , \inf_abs2_a_0[3] , \inf_abs2_5[4] , 
        \inf_abs2_a_0[4] , \inf_abs2_5[5] , \inf_abs2_a_0[5] , 
        \inf_abs2_5[10] , \inf_abs2_a_0[10] , \inf_abs2_5[13] , 
        \inf_abs2_a_0[13] , N1079, I360_un1_Y, \next_sum[17] , 
        \next_sum[0] , N_228, \state[2]_net_1 , \next_sum[1] , 
        \next_sum[2] , \next_sum[3] , \next_sum[4] , \next_sum[5] , 
        \next_sum[6] , \next_sum[7] , \next_sum[8] , \next_sum[9] , 
        \next_sum[11] , \next_sum[13] , \next_sum[14] , \next_sum[16] , 
        N1082, \next_sum[19] , N1073, \next_sum[20] , N1070, 
        \next_sum[21] , N1067, \next_sum[23] , N1061, \next_sum[24] , 
        \next_sum[25] , \next_sum[28] , \next_sum[29] , \next_sum[31] , 
        \next_sum[37] , \next_sum[38] , N282, N284, N285, N288, N290, 
        N294, N343, N293, N347, N287, N351, N278, N281, N344, N388, 
        N390, N391, I114_un1_Y, N350, N348, N346, N340, N300, N339, 
        N296, N299, N336, N315, N302, N305, N306, N308, N309, N311, 
        N349, I80_un1_Y, N353, \next_ireg_3[6] , \i_adj[0]_net_1 , 
        N722, N641, N645, N725, N648, N644, N726, N649, N729, N652, 
        N730, N653, N733, N656, N701, N694, N702, I224_un1_Y, N709, 
        N710, N717, N718, N714, N804, N807, N811, N737, N738, N815, 
        N741, N490, N493, N657, N484, N487, N795, N721, N713, N636, 
        N633, N632, N519, N523, N522_0, N520, N637, N517, N514, N617, 
        N621, N538, N541, I106_un1_Y_0, N486, N483, N640, N513_0, N516, 
        N628, I78_un1_Y, N528_0, N525_0, N529, N625, N624, N620, N537, 
        N540, N613, N616, N612, N489, N492_0, N496, N499, N495, N498_0, 
        N502, N505, N501, N504_0, N507_0, N508, N510, N511, N638, N639, 
        N642, N643, N647, N650, N651, N654, N655, N658, N480, N481, 
        N716, N635, N719, N720, N723, N646, N724, N727, N728, N731, 
        N732, N735, N736, I186_un1_Y, N662, N739, N704, N712, 
        I242_un1_Y, N801, N802, N806, N809, N810, I254_un1_Y, N813, 
        N631, N526, N711, N634, N630, N531_0, N532, N534, N535, N543, 
        N544, N546, N547, N604, N605, N618, N619, N622, N623, 
        I74_un1_Y, I76_un1_Y, N626, N627, N603, N607, N608, N609, N688, 
        N611, N690, N614, N610, N692, N615, N695, N696, N697, 
        I146_un1_Y, N699, N700, N707, N708, N715, I214_un1_Y, 
        I218_un1_Y, N703, N705, N797, N803, N805, N808, I116_un1_Y, 
        N869, I304_un1_Y, N875, I320_un1_Y, N871, \inf_abs2_5[9] , 
        \inf_abs2_a_0[9] , \inf_abs2_5[12] , \inf_abs2_a_0[12] , 
        \inf_abs2_5[15] , \inf_abs2_a_0[15] , \inf_abs2_5[16] , 
        \inf_abs2_a_0[16] , \inf_abs2_5[19] , \inf_abs2_a_0[19] , 
        \inf_abs2_5[21] , \inf_abs2_a_0[21] , \ireg[6]_net_1 , 
        \ireg[7]_net_1 , \ireg[8]_net_1 , \ireg[9]_net_1 , 
        \ireg[10]_net_1 , \ireg[11]_net_1 , \ireg[12]_net_1 , 
        \ireg[13]_net_1 , \ireg[14]_net_1 , \ireg[15]_net_1 , 
        \ireg[16]_net_1 , \ireg[25]_net_1 , \state_ns[0] , 
        \ireg[18]_net_1 , \inf_abs2_5[6] , \inf_abs2_a_0[6] , 
        \inf_abs2_5[17] , \inf_abs2_a_0[17] , \inf_abs2_5[11] , 
        \inf_abs2_a_0[11] , \inf_abs2_5[14] , \inf_abs2_a_0[14] , 
        \next_sum[33] , \next_sum[26] , N606, N660, N664, I184_un1_Y, 
        N471, N768, I156_un1_Y, N629, \next_sum[32] , \next_sum[12] , 
        N1064, \next_sum[22] , \inf_abs1_5[10] , \inf_abs1_a_2[10] , 
        \inf_abs1_5[8] , \inf_abs1_a_2[8] , \inf_abs1_5[7] , 
        \inf_abs1_a_2[7] , \inf_abs1_5[5] , \inf_abs1_a_2[5] , 
        \next_sum[15] , \next_sum[36] , \next_sum[30] , N602, N762, 
        \next_sum[35] , N550, I150_un1_Y, \next_sum[34] , 
        \next_sum[27] , \next_sum[10] , \inf_abs2_5[18] , 
        \inf_abs2_a_0[18] , \inf_abs2_5[2] , \inf_abs2_a_0[2] , 
        \inf_abs2_5[1] , \inf_abs2_a_0[1] , \inf_abs2_5[20] , 
        \inf_abs2_a_0[20] , \inf_abs2_5[8] , \inf_abs2_a_0[8] , 
        \inf_abs2_5[7] , \inf_abs2_a_0[7] , \inf_abs2_5[0] , N275, 
        N279, N357, N269, I115_un1_Y, N392, I54_un1_Y, N276, N356, 
        N355, N352, N272, \p_adj[0]_net_1 , \p_adj[1]_net_1 , 
        \p_adj[2]_net_1 , \p_adj[3]_net_1 , \p_adj[4]_net_1 , 
        \p_adj[5]_net_1 , \p_adj[6]_net_1 , \p_adj[7]_net_1 , 
        \p_adj[8]_net_1 , \p_adj[9]_net_1 , \p_adj[10]_net_1 , 
        \p_adj[11]_net_1 , \p_adj[12]_net_1 , N_6, \DWACT_FINC_E[28] , 
        \DWACT_FINC_E[13] , \DWACT_FINC_E[15] , N_7, 
        \DWACT_FINC_E[14] , N_8, \DWACT_FINC_E[9] , \DWACT_FINC_E[12] , 
        N_9_0, \DWACT_FINC_E[10] , \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[5] , N_10_0, \DWACT_FINC_E[11] , N_11_0, N_12_0, 
        N_13, \DWACT_FINC_E[8] , N_14, N_16, N_17, \DWACT_FINC_E[3] , 
        N_19, N_20, N_21, \DWACT_FINC_E[1] , N_22, N_24, N_3, 
        \DWACT_FINC_E_0[2] , \DWACT_FINC_E_0[5] , N_4, 
        \DWACT_FINC_E_0[3] , N_6_0, N_7_0, N_8_0, \DWACT_FINC_E_0[1] , 
        N_9_1, N_11_1, GND, VCC;
    
    DFN1E1C0 \sumreg[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(sum_39));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I77_Y (.A(N529), .B(N532), .Y(
        N627));
    NOR3B \preg_RNI1D2P[6]  (.A(sr_new_0_0), .B(\state[5]_net_1 ), .C(
        \preg[6]_net_1 ), .Y(\un24_next_sum_m[6] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_o3_0 (.A(
        ADD_22x22_fast_I142_Y_0_a3_3_0), .B(N513), .C(
        ADD_22x22_fast_I142_Y_0_o3_0_0), .Y(N_11));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I19_G0N (.A(\un1_next_sum[19] )
        , .B(sum_19), .Y(N528_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I14_P0N (.A(
        \un1_next_sum_iv_1[14] ), .B(\un1_next_sum_iv_2[14] ), .C(
        sum_14), .Y(N514));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I46_Y (.A(\sumreg[34]_net_1 ), 
        .B(\sumreg[35]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N596)
        );
    XA1B \sumreg_RNO[10]  (.A(N1100), .B(ADD_40x40_fast_I428_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[10] ));
    NOR3B \ireg_RNIQCJQ[10]  (.A(\state[3]_net_1 ), .B(
        \ireg[10]_net_1 ), .C(integral_1_0), .Y(\ireg_m[10] ));
    MX2 \p_adj_RNO[2]  (.A(sr_new[2]), .B(\inf_abs1_a_2[2] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[2] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I336_un1_Y (.A(N844), .B(N875), 
        .Y(I336_un1_Y));
    XA1B \sumreg_RNO[11]  (.A(N1097), .B(ADD_40x40_fast_I429_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[11] ));
    NOR3B \ireg_RNI0JJQ[16]  (.A(\state[3]_net_1 ), .B(
        \ireg[16]_net_1 ), .C(integral_1_0), .Y(\ireg_m[16] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_0 (.A(N333), .B(N330), .C(
        N329), .Y(ADD_22x22_fast_I144_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I241_Y (.A(N726), .B(N718), .Y(
        N800));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I114_Y (.A(N471), .B(
        \un1_next_sum[0] ), .C(sum_1_d0), .Y(N664));
    DFN1E1C0 \i_adj[19]  (.D(\inf_abs2_5[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[19]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I113_Y (.A(N389), .B(N396), .C(
        N388), .Y(N525));
    DFN1E1C0 \sumreg[23]  (.D(\next_sum[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_23));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I128_un1_Y_0 (.A(N383), .B(N375)
        , .Y(ADD_22x22_fast_I128_un1_Y_0));
    NOR3B inf_abs1_a_2_I_19 (.A(\DWACT_FINC_E_0[2] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[6]), .Y(N_7_0));
    OR3 \preg_RNIRS6S1[9]  (.A(\un24_next_sum_m[9] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[9] ), .Y(
        \un1_next_sum_iv_2[9] ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I33_Y (.A(\i_adj[12]_net_1 ), .B(
        \i_adj[14]_net_1 ), .C(N300), .Y(N338));
    OR2 \preg_RNIGRL33[9]  (.A(\un1_next_sum_iv_2[9] ), .B(
        \un1_next_sum_iv_1[9] ), .Y(\un1_next_sum[9] ));
    AND3 inf_abs2_a_0_I_30 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E_0[6] ));
    OR3 \ireg_RNIJK171[24]  (.A(next_sum_0_sqmuxa_2), .B(
        next_sum_0_sqmuxa_1), .C(\un1_next_sum_iv_0[24] ), .Y(
        \un1_next_sum[24] ));
    MX2 \i_adj_RNO[5]  (.A(integral[11]), .B(\inf_abs2_a_0[5] ), .S(
        integral[25]), .Y(\inf_abs2_5[5] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I304_Y (.A(I304_un1_Y), .B(N791), 
        .Y(N875));
    DFN1E1C0 \sumreg[38]  (.D(\next_sum[38] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(\sumreg[38]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I126_un1_Y_0 (.A(N371), .B(N379)
        , .Y(ADD_22x22_fast_I126_un1_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I361_Y (.A(N884), .B(
        \un1_next_sum[0] ), .C(N883), .Y(N1082));
    DFN1E1C0 \sumreg[5]  (.D(\next_sum[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNI172K[6]_net_1 ), .Q(sum_5));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I248_Y (.A(N733), .B(N726), .C(
        N725), .Y(N807));
    DFN1E1C0 \sumreg[20]  (.D(\next_sum[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_20));
    AO1 next_ireg_3_0_ADD_22x22_fast_I128_Y (.A(
        ADD_22x22_fast_I128_un1_Y_0), .B(N528), .C(
        ADD_22x22_fast_I128_Y_0), .Y(N504));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I150_un1_Y (.A(N626), .B(N623), 
        .Y(I150_un1_Y));
    NOR2 inf_abs2_a_0_I_57 (.A(integral[24]), .B(integral[25]), .Y(
        \DWACT_FINC_E[14] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I347_Y_0 (.A(N787), .B(N772), .C(
        N771), .Y(ADD_40x40_fast_I347_Y_0));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I52_Y (.A(\sumreg[32]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N602)
        );
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I199_Y (.A(N599), .B(N595), .C(
        N684), .Y(N758));
    DFN1E1C0 \sumreg[13]  (.D(\next_sum[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_13));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I76_un1_Y (.A(N528_0), .B(N532)
        , .Y(I76_un1_Y));
    OR3 \state_RNIREQ01_0[3]  (.A(next_sum_1_sqmuxa_2), .B(
        next_sum_1_sqmuxa_1), .C(next_sum_1_sqmuxa), .Y(
        \un1_next_sum_1_iv[26] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I354_Y (.A(N870), .B(N817), .C(
        N869), .Y(N1061));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I214_Y (.A(I214_un1_Y), .B(N691), 
        .Y(N773));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I353_un1_Y_0 (.A(N800), .B(
        N784), .Y(ADD_40x40_fast_I353_un1_Y_0));
    DFN1E1C0 \i_adj[2]  (.D(\inf_abs2_5[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[2]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I225_Y (.A(N702), .B(N710), .Y(
        N784));
    NOR3A inf_abs1_a_2_I_13 (.A(\DWACT_FINC_E[0] ), .B(sr_new[4]), .C(
        sr_new[3]), .Y(N_9_1));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I436_Y_0 (.A(
        \un1_next_sum_iv_1[18] ), .B(\un1_next_sum_iv_2[18] ), .C(
        sum_18), .Y(ADD_40x40_fast_I436_Y_0));
    DFN1E1C0 \sumreg[27]  (.D(\next_sum[27] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[27]_net_1 ));
    DFN1E1C0 \sumreg[10]  (.D(\next_sum[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_10));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I381_Y_2 (.A(N760), .B(N775), .C(
        ADD_40x40_fast_I381_Y_1), .Y(ADD_40x40_fast_I381_Y_2));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I308_Y (.A(N811), .B(N796), .C(
        N795), .Y(N879));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I444_Y_0 (.A(
        \sumreg[26]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I444_Y_0));
    XA1B \sumreg_RNO[22]  (.A(N1064), .B(ADD_40x40_fast_I440_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[22] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I171_Y (.A(N647), .B(N643), .Y(
        N724));
    OR2 next_ireg_3_0_ADD_22x22_fast_I11_P0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(N300));
    OR3 \preg_RNILM6S1[6]  (.A(\un24_next_sum_m[6] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[6] ), .Y(
        \un1_next_sum_iv_2[6] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I443_Y_0 (.A(
        \sumreg[25]_net_1 ), .B(\un1_next_sum_0_iv[25] ), .Y(
        ADD_40x40_fast_I443_Y_0));
    AND2 inf_abs2_a_0_I_44 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E[9] ), .Y(\DWACT_FINC_E[10] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I18_P0N (.A(
        \un1_next_sum_iv_1[18] ), .B(\un1_next_sum_iv_2[18] ), .C(
        sum_18), .Y(N526));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I166_Y (.A(N642), .B(N639), .C(
        N638), .Y(N719));
    OA1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_0_0 (.A(
        \i_adj[18]_net_1 ), .B(\i_adj[20]_net_1 ), .C(N_9), .Y(
        ADD_22x22_fast_I142_Y_0_a3_0));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I168_Y (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[8]_net_1 ), .C(N522), .Y(\next_ireg_3[14] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I384_Y_1 (.A(N766), .B(N781), .C(
        ADD_40x40_fast_I384_Y_0), .Y(ADD_40x40_fast_I384_Y_1));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I10_G0N (.A(
        \un1_next_sum_iv_1[10] ), .B(\un1_next_sum_iv_2[10] ), .C(
        sum_10), .Y(N501));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I274_un1_Y (.A(N762), .B(N777), 
        .Y(I274_un1_Y));
    XNOR2 inf_abs1_a_2_I_28 (.A(sr_new[10]), .B(N_4), .Y(
        \inf_abs1_a_2[10] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I18_G0N (.A(
        \un1_next_sum_iv_1[18] ), .B(\un1_next_sum_iv_2[18] ), .C(
        sum_18), .Y(N525_0));
    DFN1E1C0 \p_adj[4]  (.D(\inf_abs1_5[4] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[4]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_2 (.A(
        ADD_22x22_fast_I144_un1_Y_0), .B(N425), .C(
        ADD_22x22_fast_I144_Y_1), .Y(ADD_22x22_fast_I144_Y_2));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I358_Y (.A(N878), .B(N743), .C(
        N877), .Y(N1073));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I7_G0N (.A(\i_adj[7]_net_1 ), 
        .B(\i_adj[9]_net_1 ), .Y(N287));
    XNOR2 inf_abs2_a_0_I_20 (.A(integral[13]), .B(N_20), .Y(
        \inf_abs2_a_0[7] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I424_Y_0 (.A(sum_6), .B(
        \un1_next_sum[6] ), .Y(ADD_40x40_fast_I424_Y_0));
    DFN1E1C0 \sumreg[17]  (.D(\next_sum[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_17));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I257_Y_1 (.A(N475), .B(N472), 
        .C(N661), .Y(ADD_40x40_fast_I257_Y_1));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I321_Y (.A(N816), .B(
        \un1_next_sum[0] ), .C(N815), .Y(N1106));
    DFN1C0 \state[6]  (.D(\state[2]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[6]_net_1 ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I423_Y_0 (.A(sum_5), .B(
        \un1_next_sum[5] ), .Y(ADD_40x40_fast_I423_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y (.A(
        ADD_22x22_fast_I126_un1_Y_0), .B(N522), .C(
        ADD_22x22_fast_I126_Y_1), .Y(N498));
    AND3 inf_abs1_a_2_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[5] ), .Y(
        \DWACT_FINC_E[6] ));
    DFN1E1C0 \sumreg[35]  (.D(\next_sum[35] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(\sumreg[35]_net_1 ));
    MX2 \i_adj_RNO[13]  (.A(integral[19]), .B(\inf_abs2_a_0[13] ), .S(
        integral_1_0), .Y(\inf_abs2_5[13] ));
    DFN1E1C0 \sumreg[4]  (.D(\next_sum[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNI172K[6]_net_1 ), .Q(sum_4));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I166_Y_0 (.A(\i_adj[6]_net_1 ), 
        .B(\i_adj[8]_net_1 ), .Y(ADD_22x22_fast_I166_Y_0));
    XA1B \sumreg_RNO[38]  (.A(N1023), .B(ADD_40x40_fast_I456_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[38] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I160_Y (.A(N636), .B(N633), .C(
        N632), .Y(N713));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I207_Y (.A(N684), .B(N692), .Y(
        N766));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I232_Y (.A(N717), .B(N710), .C(
        N709), .Y(N791));
    NOR2 inf_abs2_a_0_I_6 (.A(integral[6]), .B(integral[7]), .Y(N_25));
    NOR3B inf_abs2_a_0_I_45 (.A(\DWACT_FINC_E[10] ), .B(
        \DWACT_FINC_E_0[6] ), .C(integral[21]), .Y(N_11_0));
    NOR3 inf_abs1_a_2_I_29 (.A(sr_new[7]), .B(sr_new[6]), .C(sr_new[8])
        , .Y(\DWACT_FINC_E_0[5] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I252_Y (.A(N737), .B(N730), .C(
        N729), .Y(N811));
    MX2 \p_adj_RNO[1]  (.A(sr_new[1]), .B(\inf_abs1_a_2[1] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[1] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I382_un1_Y (.A(N878), .B(N743), 
        .C(N846), .Y(I382_un1_Y));
    AO1 next_ireg_3_0_ADD_22x22_fast_I30_Y (.A(N302), .B(N306), .C(
        N305), .Y(N335));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I124_un1_Y (.A(N377), .B(N369), 
        .C(N424), .Y(I124_un1_Y));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I382_Y_2 (.A(I274_un1_Y), .B(
        ADD_40x40_fast_I382_Y_0), .C(I382_un1_Y), .Y(
        ADD_40x40_fast_I382_Y_2));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I330_un1_Y (.A(N838), .B(N869), 
        .Y(I330_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I237_Y (.A(N722), .B(N714), .Y(
        N796));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I12_G0N (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[12]_net_1 ), .Y(N302));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I11_G0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(N299));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I58_Y (.A(\sumreg[28]_net_1 ), 
        .B(\sumreg[29]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N608)
        );
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I257_Y (.A(
        ADD_40x40_fast_I257_Y_1), .B(N734), .Y(N816));
    OA1 next_ireg_3_0_ADD_22x22_fast_I35_Y (.A(\i_adj[12]_net_1 ), .B(
        \i_adj[10]_net_1 ), .C(N300), .Y(N340));
    OR3 \ireg_RNIGH171[21]  (.A(next_sum_0_sqmuxa_2), .B(
        next_sum_0_sqmuxa_1), .C(\un1_next_sum_iv_0[21] ), .Y(
        \un1_next_sum[21] ));
    NOR2B un1_sumreg_0_0_ADD_m8_i_a4_0_0 (.A(sum_0_d0), .B(sum_1_d0), 
        .Y(ADD_m8_i_a4_0_0));
    DFN1E1C0 \sumreg[7]  (.D(\next_sum[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNI172K[6]_net_1 ), .Q(sum_7));
    DFN1E1C0 \ireg[12]  (.D(\next_ireg_3[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[12]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I78_un1_Y (.A(N525_0), .B(N529)
        , .Y(I78_un1_Y));
    NOR3B \preg_RNIHGHP[14]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[14]_net_1 ), .Y(\un24_next_sum_m[14] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I126_Y (.A(N602), .B(I122_un1_Y), 
        .Y(N679));
    NOR2A inf_abs2_a_0_I_11 (.A(\DWACT_FINC_E_0[0] ), .B(integral[9]), 
        .Y(N_23));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I166_Y (.A(
        ADD_22x22_fast_I166_Y_0), .B(N528), .Y(\next_ireg_3[12] ));
    OR3 \preg_RNINIEQ1[16]  (.A(\un24_next_sum_m[16] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[16] ), .Y(
        \un1_next_sum_iv_2[16] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I67_Y (.A(N547), .B(N544), .Y(
        N617));
    AO1 next_ireg_3_0_ADD_22x22_fast_I38_Y (.A(N290), .B(N294), .C(
        N293), .Y(N343));
    XNOR2 inf_abs2_a_0_I_46 (.A(integral[22]), .B(N_11_0), .Y(
        \inf_abs2_a_0[16] ));
    XOR2 inf_abs1_a_2_I_5 (.A(sr_new[0]), .B(sr_new[1]), .Y(
        \inf_abs1_a_2[1] ));
    XNOR2 inf_abs1_a_2_I_23 (.A(sr_new[8]), .B(N_6_0), .Y(
        \inf_abs1_a_2[8] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I310_Y (.A(N813), .B(N798), .C(
        N797), .Y(N881));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I169_Y (.A(N641), .B(N645), .Y(
        N722));
    DFN1C0 \state[2]  (.D(\state[1]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[2]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I245_Y (.A(N722), .B(N730), .Y(
        N804));
    DFN1E1C0 \i_adj[15]  (.D(\inf_abs2_5[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[15]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I349_Y_0 (.A(N791), .B(N776), .C(
        N775), .Y(ADD_40x40_fast_I349_Y_0));
    OA1 next_ireg_3_0_ADD_22x22_fast_I41_Y (.A(\i_adj[8]_net_1 ), .B(
        \i_adj[10]_net_1 ), .C(N288), .Y(N346));
    DFN1E1C0 \i_adj[20]  (.D(\inf_abs2_5[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[20]_net_1 ));
    XNOR2 inf_abs2_a_0_I_37 (.A(integral[19]), .B(N_14), .Y(
        \inf_abs2_a_0[13] ));
    MX2 \i_adj_RNO[12]  (.A(integral[18]), .B(\inf_abs2_a_0[12] ), .S(
        integral_1_0), .Y(\inf_abs2_5[12] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I348_Y_0 (.A(N789), .B(N774), .C(
        N773), .Y(ADD_40x40_fast_I348_Y_0));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I53_Y (.A(\sumreg[31]_net_1 ), 
        .B(\sumreg[32]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N603)
        );
    AO1 next_ireg_3_0_ADD_22x22_fast_I86_Y (.A(N356), .B(N359), .C(
        N355), .Y(N394));
    AX1D next_ireg_3_0_ADD_22x22_fast_I170_Y (.A(N422), .B(I132_un1_Y), 
        .C(ADD_22x22_fast_I170_Y_0), .Y(\next_ireg_3[16] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I379_un1_Y (.A(N840), .B(N872), 
        .C(N819), .Y(I379_un1_Y));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_1 (.A(N369), .B(N376), .C(
        ADD_22x22_fast_I144_Y_0), .Y(ADD_22x22_fast_I144_Y_1));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I4_P0N (.A(\un1_next_sum[4] ), 
        .B(sum_4), .Y(N484));
    NOR2A \state_RNI5HFA_0[4]  (.A(\state[4]_net_1 ), .B(derivative_0), 
        .Y(next_sum_1_sqmuxa_1));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I213_Y (.A(N690), .B(N698), .Y(
        N772));
    DFN1E1C0 \p_adj[10]  (.D(\inf_abs1_5[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[10]_net_1 ));
    DFN1E1C0 \p_adj[5]  (.D(\inf_abs1_5[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[5]_net_1 ));
    NOR3B \ireg_RNIDA3J[15]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[15]_net_1 ), .Y(\un3_next_sum_m[15] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I164_Y (.A(N640), .B(N637), .C(
        N636), .Y(N717));
    DFN1E1C0 \sumreg[36]  (.D(\next_sum[36] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(\sumreg[36]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I56_Y (.A(\sumreg[29]_net_1 ), 
        .B(\sumreg[30]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N606)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I172_Y (.A(N648), .B(N645), .C(
        N644), .Y(N725));
    NOR2B \p_adj_RNO[12]  (.A(\inf_abs1_a_2[12] ), .B(sr_new[12]), .Y(
        \inf_abs1_5[12] ));
    OR3 \preg_RNIRMEQ1[18]  (.A(\un24_next_sum_m[18] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[18] ), .Y(
        \un1_next_sum_iv_2[18] ));
    OR3 \ireg_RNI1O151[4]  (.A(next_sum_0_sqmuxa_2), .B(
        next_sum_0_sqmuxa_1), .C(\un1_next_sum_iv_0[4] ), .Y(
        \un1_next_sum[4] ));
    NOR2B \state_RNIK76G[0]  (.A(sum_enable), .B(sum_rdy), .Y(
        \state_RNIK76G[0]_net_1 ));
    DFN1E1C0 \p_adj[0]  (.D(\inf_abs1_5[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[0]_net_1 ));
    NOR3B \preg_RNIC8BL[10]  (.A(sr_new_0_0), .B(\state[5]_net_1 ), .C(
        \preg[10]_net_1 ), .Y(\un24_next_sum_m[10] ));
    AND3 inf_abs2_a_0_I_51 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[28] ));
    DFN1E1C0 \sumreg[9]  (.D(\next_sum[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNI172K[6]_net_1 ), .Q(sum_9));
    NOR3B \preg_RNI4G2P[9]  (.A(sr_new_0_0), .B(\state[5]_net_1 ), .C(
        \preg[9]_net_1 ), .Y(\un24_next_sum_m[9] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I181_Y (.A(N657), .B(N653), .Y(
        N734));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I216_Y (.A(N701), .B(N694), .C(
        N693), .Y(N775));
    NOR3B \preg_RNI3F2P[8]  (.A(sr_new_0_0), .B(\state[5]_net_1 ), .C(
        \preg[8]_net_1 ), .Y(\un24_next_sum_m[8] ));
    OA1 un1_sumreg_0_0_ADD_m8_i_a4 (.A(N_232), .B(ADD_m8_i_o4_1), .C(
        next_sum_0_sqmuxa), .Y(ADD_m8_i_a4_4));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I4_G0N (.A(\un1_next_sum[4] ), 
        .B(sum_4), .Y(N483));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I317_Y (.A(N808), .B(N823), .C(
        N807), .Y(N1094));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I129_Y (.A(N601), .B(N605), .Y(
        N682));
    AO1 next_ireg_3_0_ADD_22x22_fast_I50_Y (.A(N272), .B(N276), .C(
        N275), .Y(N355));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I144_un1_Y_0 (.A(N377), .B(N369)
        , .C(N266), .Y(ADD_22x22_fast_I144_un1_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I34_Y (.A(N296), .B(N300), .C(
        N299), .Y(N339));
    DFN1E1C0 \sumreg[31]  (.D(\next_sum[31] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(\sumreg[31]_net_1 ));
    DFN1E1C0 \sumreg[2]  (.D(\next_sum[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNI172K[6]_net_1 ), .Q(sum_2_d0));
    DFN1E1C0 \i_adj[7]  (.D(\inf_abs2_5[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[7]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I383_Y (.A(N848), .B(N879), .C(
        ADD_40x40_fast_I383_Y_2), .Y(N1031));
    MX2 \i_adj_RNO[8]  (.A(integral[14]), .B(\inf_abs2_a_0[8] ), .S(
        integral[25]), .Y(\inf_abs2_5[8] ));
    NOR3B \preg_RNI2E2P[7]  (.A(sr_new_0_0), .B(\state[5]_net_1 ), .C(
        \preg[7]_net_1 ), .Y(\un24_next_sum_m[7] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I9_P0N (.A(\un1_next_sum[9] ), 
        .B(sum_9), .Y(N499));
    NOR3A inf_abs2_a_0_I_27 (.A(\DWACT_FINC_E_0[4] ), .B(integral[14]), 
        .C(integral[15]), .Y(N_17));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I105_Y (.A(N487), .B(N490), .Y(
        N655));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I10_G0N (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[12]_net_1 ), .Y(N296));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I351_un1_Y_0 (.A(N706), .B(
        N698), .C(N796), .Y(ADD_40x40_fast_I351_un1_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I108_Y (.A(N390), .B(N383), .C(
        N382), .Y(N422));
    MX2 \p_adj_RNO[3]  (.A(sr_new[3]), .B(\inf_abs1_a_2[3] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[3] ));
    OR3 \state_RNIF2M51[4]  (.A(next_sum_0_sqmuxa_2), .B(
        next_sum_0_sqmuxa_1), .C(N_232), .Y(N_228));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I435_Y_0 (.A(
        \un1_next_sum_iv_1[17] ), .B(\un1_next_sum_iv_2[17] ), .C(
        sum_17), .Y(ADD_40x40_fast_I435_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I146_Y (.A(I146_un1_Y), .B(N618), 
        .Y(N699));
    AND3 inf_abs2_a_0_I_48 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[11] ), .Y(N_10_0));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I197_Y_0 (.A(\sumreg[36]_net_1 )
        , .B(\sumreg[37]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(
        ADD_40x40_fast_I197_Y_0));
    DFN1E1C0 \preg[16]  (.D(\p_adj[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[16]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I135_Y (.A(N611), .B(N607), .Y(
        N688));
    DFN1E1C0 \preg[17]  (.D(\p_adj[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[17]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I9_G0N (.A(\i_adj[11]_net_1 ), 
        .B(\i_adj[9]_net_1 ), .Y(N293));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I155_Y (.A(N627), .B(N631), .Y(
        N708));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I122_un1_Y (.A(N375), .B(N367), 
        .C(N422), .Y(I122_un1_Y_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I5_P0N (.A(\i_adj[5]_net_1 ), .B(
        \i_adj[7]_net_1 ), .Y(N282));
    DFN1E1C0 \i_adj[8]  (.D(\inf_abs2_5[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[8]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I94_Y (.A(N501), .B(N505), .C(
        N504_0), .Y(N644));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I73_Y (.A(N346), .B(N342), .Y(
        N381));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I174_Y (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .C(N504), .Y(\next_ireg_3[20] ));
    DFN1E1C0 \i_adj[17]  (.D(\inf_abs2_5[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[17]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I214_un1_Y (.A(N699), .B(N692), 
        .Y(I214_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I140_Y (.A(N616), .B(N613), .C(
        N612), .Y(N693));
    OR3 \preg_RNIPUTI1[10]  (.A(\un24_next_sum_m[10] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[10] ), .Y(
        \un1_next_sum_iv_2[10] ));
    MX2 \i_adj_RNO[3]  (.A(integral[9]), .B(\inf_abs2_a_0[3] ), .S(
        integral[25]), .Y(\inf_abs2_5[3] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I74_Y (.A(I74_un1_Y), .B(N534), 
        .Y(N624));
    XNOR2 inf_abs2_a_0_I_49 (.A(integral[23]), .B(N_10_0), .Y(
        \inf_abs2_a_0[17] ));
    XNOR2 inf_abs2_a_0_I_12 (.A(integral[10]), .B(N_23), .Y(
        \inf_abs2_a_0[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I319_Y (.A(N812), .B(N745), .C(
        N811), .Y(N1100));
    XA1B \sumreg_RNO[18]  (.A(N1076), .B(ADD_40x40_fast_I436_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[18] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I383_un1_Y_0 (.A(N796), .B(
        N812), .C(N745), .Y(ADD_40x40_fast_I383_un1_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I306_Y (.A(N809), .B(N794), .C(
        N793), .Y(N877));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I224_Y (.A(I224_un1_Y), .B(N701), 
        .Y(N783));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I209_Y (.A(N686), .B(N694), .Y(
        N768));
    OR3 \ireg_RNINN071[19]  (.A(next_sum_0_sqmuxa_2), .B(
        next_sum_0_sqmuxa_1), .C(\un1_next_sum_iv_0[19] ), .Y(
        \un1_next_sum[19] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I224_un1_Y (.A(N709), .B(N702), 
        .Y(I224_un1_Y));
    NOR3B \preg_RNIIHHP[15]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[15]_net_1 ), .Y(\un24_next_sum_m[15] ));
    NOR3B \ireg_RNIVI4H[8]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[8]_net_1 ), .C(integral_0_0), .Y(\ireg_m[8] ));
    XA1 \ireg_RNISF4H[5]  (.A(integral_0_0), .B(\ireg[5]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[5] ));
    OR3 \preg_RNIR0UI1[11]  (.A(\un24_next_sum_m[11] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[11] ), .Y(
        \un1_next_sum_iv_2[11] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I383_Y_0 (.A(N681), .B(N689), .Y(
        ADD_40x40_fast_I383_Y_0));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I17_G0N (.A(
        \un1_next_sum_iv_1[17] ), .B(\un1_next_sum_iv_2[17] ), .C(
        sum_17), .Y(N522_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I356_Y (.A(N874), .B(N821), .C(
        N873), .Y(N1067));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I239_Y (.A(N716), .B(N724), .Y(
        N798));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I259_Y (.A(N738), .B(N745), .C(
        N737), .Y(N819));
    NOR3B \preg_RNIJIHP[16]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[16]_net_1 ), .Y(\un24_next_sum_m[16] ));
    NOR2B \i_adj_RNO[21]  (.A(\inf_abs2_a_0[21] ), .B(integral[25]), 
        .Y(\inf_abs2_5[21] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I116_un1_Y (.A(N472), .B(
        \un1_next_sum[0] ), .Y(I116_un1_Y));
    DFN1E1C0 \sumreg[6]  (.D(\next_sum[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNI172K[6]_net_1 ), .Q(sum_6));
    DFN1E1C0 \sumreg[0]  (.D(\next_sum[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNI172K[6]_net_1 ), .Q(sum_0_d0));
    DFN1E1C0 \preg[15]  (.D(\p_adj[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[15]_net_1 ));
    DFN1E1C0 \i_adj[10]  (.D(\inf_abs2_5[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[10]_net_1 ));
    NOR3B \ireg_RNI1HDM[18]  (.A(integral_0_0), .B(\state[3]_net_1 ), 
        .C(\ireg[18]_net_1 ), .Y(\un3_next_sum_m[18] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I452_Y_0 (.A(
        \sumreg[34]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I452_Y_0));
    DFN1E1C0 \ireg[24]  (.D(\next_ireg_3[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[24]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I271_Y (.A(N758), .B(N774), .Y(
        N842));
    XNOR2 inf_abs2_a_0_I_43 (.A(integral[21]), .B(N_12_0), .Y(
        \inf_abs2_a_0[15] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I69_Y (.A(N338), .B(N342), .Y(
        N377));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I385_Y (.A(N852), .B(N883), .C(
        ADD_40x40_fast_I385_Y_2), .Y(N1035));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I184_un1_Y (.A(N660), .B(N657), 
        .Y(I184_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I149_Y (.A(N625), .B(N621), .Y(
        N702));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I67_Y (.A(N336), .B(N340), .Y(
        N375));
    OR2 next_ireg_3_0_ADD_22x22_fast_I54_Y (.A(N269), .B(I54_un1_Y), 
        .Y(N359));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I378_Y_2 (.A(N594), .B(
        ADD_40x40_fast_I378_Y_0), .C(N679), .Y(ADD_40x40_fast_I378_Y_2)
        );
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I360_Y (.A(N881), .B(I360_un1_Y), 
        .Y(N1079));
    MX2 \p_adj_RNO[0]  (.A(sr_new[0]), .B(sr_new[0]), .S(sr_new_0_0), 
        .Y(\inf_abs1_5[0] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I384_Y_0 (.A(N691), .B(N684), .C(
        N683), .Y(ADD_40x40_fast_I384_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I182_Y (.A(N658), .B(N655), .C(
        N654), .Y(N735));
    AND3 inf_abs2_a_0_I_52 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[12] ), .Y(N_9_0));
    NOR3A inf_abs2_a_0_I_31 (.A(\DWACT_FINC_E_0[6] ), .B(integral[15]), 
        .C(integral[16]), .Y(N_16));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I163_Y (.A(N635), .B(N639), .Y(
        N716));
    AO1 next_ireg_3_0_ADD_22x22_fast_I110_Y (.A(N392), .B(N385), .C(
        N384), .Y(N424));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I197_Y (.A(N597), .B(
        ADD_40x40_fast_I197_Y_0), .C(N682), .Y(N756));
    DFN1E1C0 \i_adj[18]  (.D(\inf_abs2_5[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[18]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I91_Y (.A(N508), .B(N511), .Y(
        N641));
    OR2A un1_sumreg_0_0_ADD_40x40_fast_I25_P0N (.A(
        \un1_next_sum_0_iv[25] ), .B(\sumreg[25]_net_1 ), .Y(N547));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I144_Y (.A(N620), .B(N617), .C(
        N616), .Y(N697));
    MX2 \i_adj_RNO[16]  (.A(integral[22]), .B(\inf_abs2_a_0[16] ), .S(
        integral_1_0), .Y(\inf_abs2_5[16] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I71_Y (.A(N538), .B(N541), .Y(
        N621));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I95_Y (.A(N502), .B(N505), .Y(
        N645));
    OR2 next_ireg_3_0_ADD_22x22_fast_I13_P0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[15]_net_1 ), .Y(N306));
    OR3 \ireg_RNI2P151[5]  (.A(next_sum_0_sqmuxa_2), .B(
        next_sum_0_sqmuxa_1), .C(\un1_next_sum_iv_0[5] ), .Y(
        \un1_next_sum[5] ));
    NOR3B \ireg_RNIUH4H[7]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[7]_net_1 ), .C(integral_0_0), .Y(\ireg_m[7] ));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I161_Y (.A(\i_adj[3]_net_1 ), .B(
        \i_adj[1]_net_1 ), .C(N266), .Y(\next_ireg_3[7] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I70_Y (.A(N343), .B(N340), .C(
        N339), .Y(N378));
    NOR3B \ireg_RNIA73J[12]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[12]_net_1 ), .Y(\un3_next_sum_m[12] ));
    NOR2A \ireg_RNIG6FS_0[25]  (.A(next_sum_1_sqmuxa), .B(
        \ireg[25]_net_1 ), .Y(\un3_next_sum_m[25] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I75_Y (.A(N532), .B(N535), .Y(
        N625));
    OR3 \preg_RNI094N1[13]  (.A(\un24_next_sum_m[13] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[13] ), .Y(
        \un1_next_sum_iv_2[13] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I168_Y (.A(N644), .B(N641), .C(
        N640), .Y(N721));
    NOR3B \ireg_RNITFJQ[13]  (.A(\state[3]_net_1 ), .B(
        \ireg[13]_net_1 ), .C(integral_1_0), .Y(\ireg_m[13] ));
    MX2 \p_adj_RNO[6]  (.A(sr_new[6]), .B(\inf_abs1_a_2[6] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[6] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I379_Y_3 (.A(N756), .B(N771), .C(
        ADD_40x40_fast_I379_Y_2), .Y(ADD_40x40_fast_I379_Y_3));
    MX2 \i_adj_RNO[1]  (.A(integral[7]), .B(\inf_abs2_a_0[1] ), .S(
        integral[25]), .Y(\inf_abs2_5[1] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I75_Y (.A(N348), .B(N344), .Y(
        N383));
    GND GND_i (.Y(GND));
    OR2 next_ireg_3_0_ADD_22x22_fast_I3_P0N (.A(\i_adj[3]_net_1 ), .B(
        \i_adj[5]_net_1 ), .Y(N276));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I143_Y_0 (.A(\i_adj[17]_net_1 ), 
        .B(\i_adj[19]_net_1 ), .C(N314), .Y(ADD_22x22_fast_I143_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I348_un1_Y_0 (.A(N790), .B(
        N774), .Y(ADD_40x40_fast_I348_un1_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I244_Y (.A(N729), .B(N722), .C(
        N721), .Y(N803));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I314_Y (.A(N802), .B(N817), .C(
        N801), .Y(N1085));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I320_Y (.A(I320_un1_Y), .B(N813), 
        .Y(N1103));
    NOR3B \ireg_RNIVHJQ[15]  (.A(\state[3]_net_1 ), .B(
        \ireg[15]_net_1 ), .C(integral_1_0), .Y(\ireg_m[15] ));
    MX2 \p_adj_RNO[5]  (.A(sr_new[5]), .B(\inf_abs1_a_2[5] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[5] ));
    NOR2B \ireg_RNIG6FS[25]  (.A(\ireg[25]_net_1 ), .B(
        next_sum_0_sqmuxa), .Y(\ireg_m[25] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I378_Y_3 (.A(N754), .B(N769), .C(
        ADD_40x40_fast_I378_Y_2), .Y(ADD_40x40_fast_I378_Y_3));
    DFN1C0 \state[5]  (.D(\state[4]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[5]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I78_Y (.A(N351), .B(N348), .C(
        N347), .Y(N386));
    NOR2 inf_abs2_a_0_I_21 (.A(integral[12]), .B(integral[13]), .Y(
        \DWACT_FINC_E[3] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I418_Y_0 (.A(sum_0_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I418_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I87_Y (.A(N517), .B(N514), .Y(
        N637));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I384_Y_2 (.A(
        ADD_40x40_fast_I384_un1_Y_0), .B(N850), .C(
        ADD_40x40_fast_I384_Y_1), .Y(ADD_40x40_fast_I384_Y_2));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I29_Y (.A(N306), .B(N309), .Y(
        N334));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I22_P0N (.A(sum_22), .B(
        \un1_next_sum[22] ), .Y(N538));
    NOR3A inf_abs1_a_2_I_31 (.A(\DWACT_FINC_E[6] ), .B(sr_new[9]), .C(
        sr_new[10]), .Y(N_3));
    OA1 next_ireg_3_0_ADD_22x22_fast_I27_Y (.A(\i_adj[17]_net_1 ), .B(
        \i_adj[15]_net_1 ), .C(N309), .Y(N332));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I223_Y (.A(N700), .B(N708), .Y(
        N782));
    DFN1E1C0 \ireg[6]  (.D(\next_ireg_3[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[6]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I349_un1_Y_0 (.A(N792), .B(
        N776), .Y(ADD_40x40_fast_I349_un1_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I294_un1_Y (.A(N797), .B(N782), 
        .Y(I294_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I23_G0N (.A(\un1_next_sum[23] )
        , .B(sum_23), .Y(N540));
    DFN1E1C0 \preg[6]  (.D(\p_adj[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[6]_net_1 ));
    NOR3B \ireg_RNI0GDM[17]  (.A(integral_0_0), .B(\state[3]_net_1 ), 
        .C(\ireg[17]_net_1 ), .Y(\un3_next_sum_m[17] ));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I36_Y (.A(N293), .B(
        \i_adj[12]_net_1 ), .C(\i_adj[10]_net_1 ), .Y(N341));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I146_un1_Y (.A(N622), .B(N619), 
        .Y(I146_un1_Y));
    AO1 \preg_RNINF6D1[10]  (.A(\preg[10]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[10] ), .Y(
        \un1_next_sum_iv_1[10] ));
    NOR2 inf_abs1_a_2_I_6 (.A(sr_new[0]), .B(sr_new[1]), .Y(N_12));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I1_G0N (.A(\i_adj[1]_net_1 ), 
        .B(\i_adj[3]_net_1 ), .Y(N269));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I318_Y (.A(N810), .B(N743), .C(
        N809), .Y(N1097));
    OR2 next_ireg_3_0_ADD_22x22_fast_I114_Y (.A(I114_un1_Y), .B(N390), 
        .Y(N528));
    AO13 un1_sumreg_0_0_ADD_40x40_fast_I64_Y (.A(\sumreg[26]_net_1 ), 
        .B(N546), .C(\un1_next_sum_1_iv[26] ), .Y(N614));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I457_Y_0 (.A(sum_39), .B(
        \un1_next_sum_1_iv[26] ), .Y(ADD_40x40_fast_I457_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I186_un1_Y (.A(N662), .B(N659), 
        .Y(I186_un1_Y));
    XA1B \sumreg_RNO[34]  (.A(N1031), .B(ADD_40x40_fast_I452_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[34] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I81_Y (.A(N354), .B(N350), .Y(
        N389));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I128_Y (.A(N604), .B(N600), .Y(
        N681));
    OR3 \state_RNIREQ01[3]  (.A(next_sum_1_sqmuxa_2), .B(
        next_sum_1_sqmuxa_1), .C(next_sum_1_sqmuxa), .Y(
        \un1_next_sum_1_iv_0[26] ));
    DFN1E1C0 \sumreg[29]  (.D(\next_sum[29] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[29]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I99_Y (.A(N496), .B(N499), .Y(
        N649));
    NOR3B \preg_RNIKJHP[17]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[17]_net_1 ), .Y(\un24_next_sum_m[17] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I169_Y_0 (.A(\i_adj[9]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(ADD_22x22_fast_I169_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I226_Y (.A(N711), .B(N704), .C(
        N703), .Y(N785));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I442_Y_0 (.A(\sumreg[24]_net_1 )
        , .B(\un1_next_sum[24] ), .Y(ADD_40x40_fast_I442_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I212_Y (.A(N697), .B(N690), .C(
        N689), .Y(N771));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I79_Y (.A(N529), .B(N526), .Y(
        N629));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I167_Y (.A(N643), .B(N639), .Y(
        N720));
    NOR3 inf_abs1_a_2_I_10 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2])
        , .Y(\DWACT_FINC_E[0] ));
    DFN1C0 \state_0[3]  (.D(\state[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_0[3]_net_1 ));
    DFN1E1C0 \ireg[21]  (.D(\next_ireg_3[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[21]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I281_Y (.A(N768), .B(N784), .Y(
        N852));
    OR3 \preg_RNIPQ6S1[8]  (.A(\un24_next_sum_m[8] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[8] ), .Y(
        \un1_next_sum_iv_2[8] ));
    XNOR2 inf_abs2_a_0_I_32 (.A(integral[17]), .B(N_16), .Y(
        \inf_abs2_a_0[11] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I350_un1_Y_0 (.A(N794), .B(
        N778), .Y(ADD_40x40_fast_I350_un1_Y_0));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I430_Y_0 (.A(
        \un1_next_sum_iv_1[12] ), .B(\un1_next_sum_iv_2[12] ), .C(
        sum_12), .Y(ADD_40x40_fast_I430_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I217_Y (.A(N694), .B(N702), .Y(
        N776));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I378_un1_Y (.A(N817), .B(N870), 
        .C(N838), .Y(I378_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I275_Y (.A(N762), .B(N778), .Y(
        N846));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I15_P0N (.A(
        \un1_next_sum_iv_1[15] ), .B(\un1_next_sum_iv_2[15] ), .C(
        sum_15), .Y(N517));
    XA1B \sumreg_RNO[27]  (.A(N1049), .B(ADD_40x40_fast_I445_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[27] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I74_Y (.A(N347), .B(N344), .C(
        N343), .Y(N382));
    DFN1E1C0 \sumreg[19]  (.D(\next_sum[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_19));
    OR3 \preg_RNIU64N1[12]  (.A(\un24_next_sum_m[12] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[12] ), .Y(
        \un1_next_sum_iv_2[12] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I422_Y_0 (.A(sum_4), .B(
        \un1_next_sum[4] ), .Y(ADD_40x40_fast_I422_Y_0));
    NOR3B \preg_RNID9BL[11]  (.A(sr_new_0_0), .B(\state[5]_net_1 ), .C(
        \preg[11]_net_1 ), .Y(\un24_next_sum_m[11] ));
    DFN1E1C0 \sumreg[8]  (.D(\next_sum[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNI172K[6]_net_1 ), .Q(sum_8));
    DFN1E1C0 \sumreg[28]  (.D(\next_sum[28] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[28]_net_1 ));
    XA1 \ireg_RNIDB4J[24]  (.A(integral_0_0), .B(\ireg[24]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[24] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I304_un1_Y (.A(N807), .B(N792), 
        .Y(I304_un1_Y));
    XA1B \sumreg_RNO[0]  (.A(N_228), .B(ADD_40x40_fast_I418_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[0] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I451_Y_0 (.A(
        \sumreg[33]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I451_Y_0));
    OR3 un1_sumreg_0_0_ADD_m8_i_1 (.A(next_sum_0_sqmuxa_2), .B(
        next_sum_0_sqmuxa_1), .C(ADD_m8_i_a4_0_1), .Y(ADD_m8_i_1));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I143_Y (.A(N615), .B(N619), .Y(
        N696));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_1_0 (.A(
        ADD_22x22_fast_I142_Y_0_a3_0), .B(N330), .Y(
        ADD_22x22_fast_I142_Y_0_a3_1));
    XA1 \ireg_RNIRE4H[4]  (.A(integral_0_0), .B(\ireg[4]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[4] ));
    DFN1C0 \state_2[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_2[2]_net_1 ));
    DFN1E1C0 \sumreg[18]  (.D(\next_sum[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_18));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I380_Y_1 (.A(I122_un1_Y), .B(
        N594), .C(N683), .Y(ADD_40x40_fast_I380_Y_1));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I61_Y (.A(\sumreg[28]_net_1 ), 
        .B(\sumreg[27]_net_1 ), .C(\un1_next_sum_1_iv[26] ), .Y(N611));
    NOR3B \ireg_RNI0K4H[9]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[9]_net_1 ), .C(integral_0_0), .Y(\ireg_m[9] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I6_G0N (.A(\i_adj[8]_net_1 ), 
        .B(\i_adj[6]_net_1 ), .Y(N284));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I162_Y (.A(\i_adj[4]_net_1 ), .B(
        \i_adj[2]_net_1 ), .C(N359), .Y(\next_ireg_3[8] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I21_P0N (.A(\un1_next_sum[21] ), 
        .B(sum_21), .Y(N535));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I243_Y (.A(N720), .B(N728), .Y(
        N802));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I127_Y (.A(N599), .B(N603), .Y(
        N680));
    DFN1E1C0 \p_adj[3]  (.D(\inf_abs1_5[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[3]_net_1 ));
    DFN1E1C0 \ireg[10]  (.D(\next_ireg_3[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[10]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I49_Y (.A(N276), .B(N279), .Y(
        N354));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I65_Y (.A(N550), .B(N547), .Y(
        N615));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I47_Y (.A(N279), .B(N282), .Y(
        N352));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I101_Y (.A(N496), .B(N493), .Y(
        N651));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I12_P0N (.A(
        \un1_next_sum_iv_1[12] ), .B(\un1_next_sum_iv_2[12] ), .C(
        sum_12), .Y(N508));
    AND3 inf_abs2_a_0_I_22 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_19));
    DFN1E1C0 \sumreg[1]  (.D(\next_sum[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNI172K[6]_net_1 ), .Q(sum_1_d0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I449_Y_0 (.A(
        \sumreg[31]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I449_Y_0));
    XA1B \sumreg_RNO[20]  (.A(N1070), .B(ADD_40x40_fast_I438_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[20] ));
    DFN1E1C0 \sumreg_0[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(sum_0_0));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I47_Y (.A(\sumreg[35]_net_1 ), 
        .B(\sumreg[34]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N597)
        );
    XNOR2 inf_abs1_a_2_I_32 (.A(sr_new[11]), .B(N_3), .Y(
        \inf_abs1_a_2[11] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I187_Y_0 (.A(\un1_next_sum[0] ), 
        .B(sum_2_d0), .C(N475), .Y(ADD_40x40_fast_I187_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I148_Y (.A(N624), .B(N621), .C(
        N620), .Y(N701));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I165_Y (.A(
        ADD_22x22_fast_I165_Y_0), .B(N531), .Y(\next_ireg_3[11] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I13_G0N (.A(
        \un1_next_sum_iv_1[13] ), .B(\un1_next_sum_iv_2[13] ), .C(
        sum_13), .Y(N510));
    XA1B \sumreg_RNO[21]  (.A(N1067), .B(ADD_40x40_fast_I439_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[21] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_3_0 (.A(N338), .B(
        N334), .Y(ADD_22x22_fast_I142_Y_0_a3_3_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I131_Y (.A(N603), .B(N607), .Y(
        N684));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I303_Y (.A(N806), .B(N790), .Y(
        N874));
    XNOR2 inf_abs1_a_2_I_20 (.A(sr_new[7]), .B(N_7_0), .Y(
        \inf_abs1_a_2[7] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I438_Y_0 (.A(sum_20), .B(
        \un1_next_sum[20] ), .Y(ADD_40x40_fast_I438_Y_0));
    DFN1E1C0 \sumreg[25]  (.D(\next_sum[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[25]_net_1 ));
    AO1 \preg_RNITL6D1[13]  (.A(\preg[13]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[13] ), .Y(
        \un1_next_sum_iv_1[13] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I246_Y (.A(N731), .B(N724), .C(
        N723), .Y(N805));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I151_Y (.A(N623), .B(N627), .Y(
        N704));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I176_Y (.A(N652), .B(N649), .C(
        N648), .Y(N729));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I347_Y (.A(
        ADD_40x40_fast_I347_un1_Y_0), .B(N1088), .C(
        ADD_40x40_fast_I347_Y_0), .Y(N1040));
    DFN1E1C0 \ireg[23]  (.D(\next_ireg_3[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[23]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I106_un1_Y (.A(N381), .B(N388), 
        .Y(I106_un1_Y));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I429_Y_0 (.A(
        \un1_next_sum_iv_1[11] ), .B(\un1_next_sum_iv_2[11] ), .C(
        sum_11), .Y(ADD_40x40_fast_I429_Y_0));
    OR2 un1_sumreg_0_0_ADD_m8_i (.A(ADD_m8_i_1), .B(ADD_m8_i_a4_4), .Y(
        N743));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I9_G0N (.A(\un1_next_sum[9] ), 
        .B(sum_9), .Y(N498_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I447_Y_0 (.A(
        \sumreg[29]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I447_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I353_Y (.A(
        ADD_40x40_fast_I353_un1_Y_0), .B(N1106), .C(
        ADD_40x40_fast_I353_Y_0), .Y(N1058));
    AND3 inf_abs2_a_0_I_60 (.A(integral_i[24]), .B(integral_i[25]), .C(
        integral_i[25]), .Y(\DWACT_FINC_E[15] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I170_Y (.A(N646), .B(N643), .C(
        N642), .Y(N723));
    DFN1E1C0 \sumreg[15]  (.D(\next_sum[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_15));
    DFN1E1C0 \ireg[5]  (.D(\i_adj[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[5]_net_1 ));
    DFN1E1C0 \ireg[25]  (.D(\next_ireg_3[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[25]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0 (.A(
        ADD_22x22_fast_I142_Y_0_a3_1), .B(N_11), .C(
        ADD_22x22_fast_I142_Y_0_1), .Y(N492));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I353_Y_0 (.A(N799), .B(N784), .C(
        N783), .Y(ADD_40x40_fast_I353_Y_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I16_P0N (.A(\i_adj[18]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .Y(N315));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I5_G0N (.A(\un1_next_sum[5] ), 
        .B(sum_5), .Y(N486));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I427_Y_0 (.A(sum_9), .B(
        \un1_next_sum[9] ), .Y(ADD_40x40_fast_I427_Y_0));
    DFN1E1C0 \p_adj[9]  (.D(\inf_abs1_5[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[9]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I80_un1_Y (.A(N353), .B(N350), 
        .Y(I80_un1_Y));
    XNOR2 inf_abs1_a_2_I_17 (.A(sr_new[6]), .B(N_8_0), .Y(
        \inf_abs1_a_2[6] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I163_Y (.A(
        ADD_22x22_fast_I163_Y_0), .B(N396), .Y(\next_ireg_3[9] ));
    MX2 \i_adj_RNO[14]  (.A(integral[20]), .B(\inf_abs2_a_0[14] ), .S(
        integral_1_0), .Y(\inf_abs2_5[14] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I69_Y (.A(N544), .B(N541), .Y(
        N619));
    XA1B \sumreg_RNO[14]  (.A(N1088), .B(ADD_40x40_fast_I432_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[14] ));
    XA1B \sumreg_RNO[35]  (.A(N1029), .B(ADD_40x40_fast_I453_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[35] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I349_Y (.A(
        ADD_40x40_fast_I349_un1_Y_0), .B(N1094), .C(
        ADD_40x40_fast_I349_Y_0), .Y(N1046));
    DFN1C0 \state[4]  (.D(\state_0[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[4]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I147_Y (.A(N623), .B(N619), .Y(
        N700));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I8_G0N (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[8]_net_1 ), .Y(N290));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_0 (.A(\i_adj[18]_net_1 )
        , .B(\i_adj[20]_net_1 ), .C(N_14_1), .Y(
        ADD_22x22_fast_I142_Y_0_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I9_P0N (.A(\i_adj[11]_net_1 ), .B(
        \i_adj[9]_net_1 ), .Y(N294));
    DFN1E1C0 \sumreg[26]  (.D(\next_sum[26] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[26]_net_1 ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I441_Y_0 (.A(sum_23), .B(
        \un1_next_sum[23] ), .Y(ADD_40x40_fast_I441_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I179_Y (.A(N655), .B(N651), .Y(
        N732));
    XA1B \sumreg_RNO[7]  (.A(N817), .B(ADD_40x40_fast_I425_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[7] ));
    OR3 \preg_RNINO6S1[7]  (.A(\un24_next_sum_m[7] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[7] ), .Y(
        \un1_next_sum_iv_2[7] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I11_P0N (.A(
        \un1_next_sum_iv_1[11] ), .B(\un1_next_sum_iv_2[11] ), .C(
        sum_11), .Y(N505));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I267_Y (.A(N754), .B(N770), .Y(
        N838));
    AO1 next_ireg_3_0_ADD_22x22_fast_I128_Y_0 (.A(N382), .B(N375), .C(
        N374), .Y(ADD_22x22_fast_I128_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I90_Y (.A(N507_0), .B(N511), .C(
        N510), .Y(N640));
    DFN1E1C0 \ireg[17]  (.D(\next_ireg_3[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[17]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I316_Y (.A(N806), .B(N821), .C(
        N805), .Y(N1091));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I305_Y (.A(N808), .B(N792), .Y(
        N876));
    OR3 \preg_RNI4D4N1[15]  (.A(\un24_next_sum_m[15] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[15] ), .Y(
        \un1_next_sum_iv_2[15] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I381_Y (.A(
        ADD_40x40_fast_I381_Y_2), .B(I381_un1_Y), .C(I336_un1_Y), .Y(
        N1027));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I219_Y (.A(N704), .B(N696), .Y(
        N778));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I102_Y (.A(N489), .B(N493), .C(
        N492_0), .Y(N652));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I70_Y (.A(N537), .B(N541), .C(
        N540), .Y(N620));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I21_G0N (.A(\un1_next_sum[21] )
        , .B(sum_21), .Y(N534));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I195_Y (.A(N595), .B(
        ADD_40x40_fast_I195_Y_0), .C(N680), .Y(N754));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I421_Y_0 (.A(sum_3), .B(N743), 
        .Y(ADD_40x40_fast_I421_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I174_Y (.A(N650), .B(N647), .C(
        N646), .Y(N727));
    XA1 \ireg_RNIHE3J[19]  (.A(integral_0_0), .B(\ireg[19]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[19] ));
    DFN1E1C0 \sumreg[16]  (.D(\next_sum[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_16));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I16_G0N (.A(\i_adj[18]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .Y(N314));
    XNOR2 inf_abs2_a_0_I_14 (.A(integral[11]), .B(N_22), .Y(
        \inf_abs2_a_0[5] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I355_Y (.A(N872), .B(N819), .C(
        N871), .Y(N1064));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I132_Y (.A(N608), .B(N604), .Y(
        N685));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I2_G0N (.A(\i_adj[4]_net_1 ), 
        .B(\i_adj[2]_net_1 ), .Y(N272));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I152_Y (.A(N628), .B(N625), .C(
        N624), .Y(N705));
    MX2 \p_adj_RNO[8]  (.A(sr_new[8]), .B(\inf_abs1_a_2[8] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[8] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I3_P0N (.A(sum_3), .B(
        \un1_next_sum[0] ), .Y(N481));
    AO1 next_ireg_3_0_ADD_22x22_fast_I76_Y (.A(N349), .B(N346), .C(
        N345), .Y(N384));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I352_un1_Y (.A(
        ADD_40x40_fast_I352_un1_Y_0), .B(N1103), .Y(I352_un1_Y));
    DFN1E1C0 \sumreg[21]  (.D(\next_sum[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_21));
    MX2 \p_adj_RNO[7]  (.A(sr_new[7]), .B(\inf_abs1_a_2[7] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[7] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I84_Y (.A(N516), .B(N520), .C(
        N519), .Y(N634));
    AO1 next_ireg_3_0_ADD_22x22_fast_I42_Y (.A(N284), .B(N288), .C(
        N287), .Y(N347));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I222_Y (.A(N707), .B(N700), .C(
        N699), .Y(N781));
    XA1B \sumreg_RNO[36]  (.A(N1027), .B(ADD_40x40_fast_I454_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[36] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I1_P0N (.A(sum_1_d0), .B(
        \un1_next_sum[0] ), .Y(N475));
    OA1 next_ireg_3_0_ADD_22x22_fast_I31_Y (.A(\i_adj[12]_net_1 ), .B(
        \i_adj[14]_net_1 ), .C(N306), .Y(N336));
    AO1 next_ireg_3_0_ADD_22x22_fast_I129_Y (.A(
        ADD_22x22_fast_I129_un1_Y_0), .B(N531), .C(
        ADD_22x22_fast_I129_Y_0), .Y(N507));
    NOR3 \state_RNI172K[6]  (.A(sum_rdy), .B(\state[6]_net_1 ), .C(
        \state[1]_net_1 ), .Y(\state_RNI172K[6]_net_1 ));
    DFN1E1C0 \p_adj[1]  (.D(\inf_abs1_5[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[1]_net_1 ));
    NOR3A inf_abs1_a_2_I_27 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .C(
        sr_new[9]), .Y(N_4));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I186_Y (.A(I186_un1_Y), .B(N658), 
        .Y(N739));
    NOR2 inf_abs2_a_0_I_15 (.A(integral[9]), .B(integral[10]), .Y(
        \DWACT_FINC_E[1] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I434_Y_0 (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(ADD_40x40_fast_I434_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I227_Y (.A(N704), .B(N712), .Y(
        N786));
    DFN1E1C0 \p_adj[7]  (.D(\inf_abs1_5[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[7]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I299_Y (.A(N802), .B(N786), .Y(
        N870));
    DFN1E1C0 \sumreg[11]  (.D(\next_sum[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_11));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I433_Y_0 (.A(
        \un1_next_sum_iv_1[15] ), .B(\un1_next_sum_iv_2[15] ), .C(
        sum_15), .Y(ADD_40x40_fast_I433_Y_0));
    OR3 \preg_RNI2B4N1[14]  (.A(\un24_next_sum_m[14] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[14] ), .Y(
        \un1_next_sum_iv_2[14] ));
    NOR3B \ireg_RNIUGJQ[14]  (.A(\state[3]_net_1 ), .B(
        \ireg[14]_net_1 ), .C(integral_1_0), .Y(\ireg_m[14] ));
    XA1B \sumreg_RNO[33]  (.A(N1033), .B(ADD_40x40_fast_I451_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[33] ));
    DFN1E1C0 \ireg[19]  (.D(\next_ireg_3[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[19]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I320_un1_Y (.A(N814), .B(N666), 
        .Y(I320_un1_Y));
    MX2 \i_adj_RNO[10]  (.A(integral[16]), .B(\inf_abs2_a_0[10] ), .S(
        integral_0_0), .Y(\inf_abs2_5[10] ));
    XNOR2 inf_abs2_a_0_I_40 (.A(integral[20]), .B(N_13), .Y(
        \inf_abs2_a_0[14] ));
    NOR3B \ireg_RNIGPKO[7]  (.A(integral_1_0), .B(\state[3]_net_1 ), 
        .C(\ireg[7]_net_1 ), .Y(\un3_next_sum_m[7] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I385_Y_0 (.A(N693), .B(N686), .C(
        N685), .Y(ADD_40x40_fast_I385_Y_0));
    NOR3B \ireg_RNISEJQ[12]  (.A(\state[3]_net_1 ), .B(
        \ireg[12]_net_1 ), .C(integral_1_0), .Y(\ireg_m[12] ));
    AND3 inf_abs2_a_0_I_54 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E[9] ), .C(\DWACT_FINC_E[12] ), .Y(
        \DWACT_FINC_E[13] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I180_Y (.A(N656), .B(N653), .C(
        N652), .Y(N733));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I167_Y (.A(\i_adj[7]_net_1 ), .B(
        \i_adj[9]_net_1 ), .C(N525), .Y(\next_ireg_3[13] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I57_Y (.A(\sumreg[30]_net_1 ), 
        .B(\sumreg[29]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N607)
        );
    DFN1C0 \state[1]  (.D(\state_RNIK76G[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[1]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I382_Y (.A(N846), .B(N877), .C(
        ADD_40x40_fast_I382_Y_2), .Y(N1029));
    MX2 \p_adj_RNO[10]  (.A(sr_new[10]), .B(\inf_abs1_a_2[10] ), .S(
        sr_new_1_0), .Y(\inf_abs1_5[10] ));
    DFN1E1C0 \ireg[22]  (.D(\next_ireg_3[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[22]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I20_P0N (.A(\un1_next_sum[20] ), 
        .B(sum_20), .Y(N532));
    AX1D next_ireg_3_0_ADD_22x22_fast_I169_Y (.A(N424), .B(I133_un1_Y), 
        .C(ADD_22x22_fast_I169_Y_0), .Y(\next_ireg_3[15] ));
    NOR3B \ireg_RNIB83J[13]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[13]_net_1 ), .Y(\un3_next_sum_m[13] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I114_un1_Y (.A(N391), .B(N359), 
        .Y(I114_un1_Y));
    NOR3B inf_abs2_a_0_I_16 (.A(\DWACT_FINC_E[1] ), .B(
        \DWACT_FINC_E_0[0] ), .C(integral[11]), .Y(N_21));
    NOR3B inf_abs2_a_0_I_55 (.A(\DWACT_FINC_E[13] ), .B(
        \DWACT_FINC_E[28] ), .C(integral[24]), .Y(N_8));
    DFN1E1C0 \preg[13]  (.D(\p_adj[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[13]_net_1 ));
    DFN1E1C0 \i_adj[6]  (.D(\inf_abs2_5[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[6]_net_1 ));
    DFN1E1C0 \i_adj[4]  (.D(\inf_abs2_5[4] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[4]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I63_Y (.A(N336), .B(N332), .Y(
        N371));
    NOR3C un1_sumreg_0_0_ADD_m8_i_a4_0 (.A(ADD_m8_i_a4_0_0), .B(
        sum_2_d0), .C(N_232), .Y(ADD_m8_i_a4_0_1));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I230_Y (.A(N715), .B(N708), .C(
        N707), .Y(N789));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I81_Y (.A(N523), .B(N526), .Y(
        N631));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I379_Y_2 (.A(N596), .B(
        ADD_40x40_fast_I379_Y_0), .C(N681), .Y(ADD_40x40_fast_I379_Y_2)
        );
    MX2 \i_adj_RNO[18]  (.A(integral[24]), .B(\inf_abs2_a_0[18] ), .S(
        integral_1_0), .Y(\inf_abs2_5[18] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I250_Y (.A(N735), .B(N728), .C(
        N727), .Y(N809));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I456_Y_0 (.A(
        \sumreg[38]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I456_Y_0));
    NOR2A inf_abs1_a_2_I_11 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .Y(
        N_10));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I348_Y (.A(
        ADD_40x40_fast_I348_un1_Y_0), .B(N1091), .C(
        ADD_40x40_fast_I348_Y_0), .Y(N1043));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I165_Y (.A(N641), .B(N637), .Y(
        N718));
    XA1 \ireg_RNI974J[20]  (.A(integral_0_0), .B(\ireg[20]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[20] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I381_Y_1 (.A(N596), .B(N600), .C(
        N685), .Y(ADD_40x40_fast_I381_Y_1));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I92_Y (.A(N504_0), .B(N508), .C(
        N507_0), .Y(N642));
    NOR2A \state_RNI1OD9_0[5]  (.A(\state[5]_net_1 ), .B(sr_new[12]), 
        .Y(next_sum_1_sqmuxa_2));
    DFN1E1C0 \i_adj[9]  (.D(\inf_abs2_5[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[9]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I85_Y (.A(N517), .B(N520), .Y(
        N635));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I11_G0N (.A(
        \un1_next_sum_iv_1[11] ), .B(\un1_next_sum_iv_2[11] ), .C(
        sum_11), .Y(N504_0));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I201_Y (.A(N597), .B(N601), .C(
        N686), .Y(N760));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I72_Y (.A(N534), .B(N538), .C(
        N537), .Y(N622));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I0_S (.A(\i_adj[0]_net_1 ), .B(
        \i_adj[2]_net_1 ), .Y(\next_ireg_3[6] ));
    DFN1E1C0 \i_adj[3]  (.D(\inf_abs2_5[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[3]_net_1 ));
    XA1B \sumreg_RNO[15]  (.A(N1085), .B(ADD_40x40_fast_I433_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[15] ));
    NOR3B \preg_RNILKHP[18]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[18]_net_1 ), .Y(\un24_next_sum_m[18] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I242_Y (.A(I242_un1_Y), .B(N719), 
        .Y(N801));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y_1 (.A(N371), .B(N378), .C(
        ADD_22x22_fast_I126_Y_0), .Y(ADD_22x22_fast_I126_Y_1));
    OR2 next_ireg_3_0_ADD_22x22_fast_I14_P0N (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .Y(N309));
    OA1 next_ireg_3_0_ADD_22x22_fast_I51_Y (.A(\i_adj[2]_net_1 ), .B(
        \i_adj[4]_net_1 ), .C(N276), .Y(N356));
    AX1D next_ireg_3_0_ADD_22x22_fast_I178_Y (.A(I122_un1_Y_0), .B(
        ADD_22x22_fast_I143_Y_3), .C(ADD_22x22_fast_I178_Y_0), .Y(
        \next_ireg_3[24] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I231_Y (.A(N716), .B(N708), .Y(
        N790));
    XA1B \state_RNIEDA1E9[2]  (.A(N1021), .B(ADD_40x40_fast_I457_Y_0), 
        .C(\state[2]_net_1 ), .Y(\next_sum[39] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I184_Y (.A(I184_un1_Y), .B(N656), 
        .Y(N737));
    XNOR2 inf_abs2_a_0_I_56 (.A(integral[25]), .B(N_8), .Y(
        \inf_abs2_a_0[19] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I87_Y (.A(I54_un1_Y), .B(N357), 
        .Y(N396));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I251_Y (.A(N736), .B(N728), .Y(
        N810));
    DFN1E1C0 \sumreg[34]  (.D(\next_sum[34] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(\sumreg[34]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I247_Y (.A(N724), .B(N732), .Y(
        N806));
    DFN1C0 \state_0[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_0[2]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I60_Y (.A(\sumreg[27]_net_1 ), 
        .B(\sumreg[28]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N610)
        );
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I385_un1_Y (.A(N884), .B(
        \un1_next_sum[0] ), .C(N852), .Y(I385_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I173_Y (.A(N645), .B(N649), .Y(
        N726));
    OR2 next_ireg_3_0_ADD_22x22_fast_I6_P0N (.A(\i_adj[8]_net_1 ), .B(
        \i_adj[6]_net_1 ), .Y(N285));
    DFN1E1C0 \ireg[7]  (.D(\next_ireg_3[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[7]_net_1 ));
    XA1B \sumreg_RNO[28]  (.A(N1046), .B(ADD_40x40_fast_I446_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[28] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I380_un1_Y (.A(N821), .B(N874), 
        .C(N842), .Y(I380_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I238_Y (.A(N723), .B(N716), .C(
        N715), .Y(N797));
    XA1B \sumreg_RNO[3]  (.A(\un1_next_sum[0] ), .B(
        ADD_40x40_fast_I421_Y_0), .C(\state[2]_net_1 ), .Y(
        \next_sum[3] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I269_Y (.A(N756), .B(N772), .Y(
        N840));
    DFN1E1C0 \preg[7]  (.D(\p_adj[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[7]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I44_Y (.A(\sumreg[35]_net_1 ), 
        .B(\sumreg[36]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N594)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I258_Y (.A(N736), .B(N743), .C(
        N735), .Y(N817));
    OR3 next_ireg_3_0_ADD_22x22_fast_I131_Y (.A(I131_un1_Y), .B(
        ADD_22x22_fast_I131_Y_0), .C(I106_un1_Y), .Y(N513));
    DFN1E1C0 \ireg[16]  (.D(\next_ireg_3[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[16]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I273_Y (.A(N760), .B(N776), .Y(
        N844));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I195_Y_0 (.A(\sumreg[37]_net_1 )
        , .B(\sumreg[38]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(
        ADD_40x40_fast_I195_Y_0));
    XA1B \sumreg_RNO[32]  (.A(N1035), .B(ADD_40x40_fast_I450_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[32] ));
    DFN1E1C0 \preg[10]  (.D(\p_adj[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[10]_net_1 ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I163_Y_0 (.A(\i_adj[5]_net_1 ), 
        .B(\i_adj[3]_net_1 ), .Y(ADD_22x22_fast_I163_Y_0));
    DFN1E1C0 \preg[18]  (.D(\p_adj[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[18]_net_1 ));
    AO1 \preg_RNIRJ6D1[12]  (.A(\preg[12]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[12] ), .Y(
        \un1_next_sum_iv_1[12] ));
    NOR3 inf_abs2_a_0_I_18 (.A(integral[10]), .B(integral[9]), .C(
        integral[11]), .Y(\DWACT_FINC_E[2] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I6_P0N (.A(\un1_next_sum[6] ), 
        .B(sum_6), .Y(N490));
    XA1B \sumreg_RNO[8]  (.A(N1106), .B(ADD_40x40_fast_I426_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[8] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I23_Y (.A(N315), .B(N_9), .Y(
        N328));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I384_un1_Y_0 (.A(N798), .B(
        N814), .C(N666), .Y(ADD_40x40_fast_I384_un1_Y_0));
    OR3 \state_RNIREQ01_1[3]  (.A(next_sum_0_sqmuxa_2), .B(
        next_sum_0_sqmuxa_1), .C(next_sum_0_sqmuxa), .Y(
        \un1_next_sum[0] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I178_Y (.A(N654), .B(N651), .C(
        N650), .Y(N731));
    NOR2B inf_abs2_a_0_I_34 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .Y(N_15));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I98_Y (.A(N495), .B(N499), .C(
        N498_0), .Y(N648));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I7_P0N (.A(
        \un1_next_sum_iv_1[7] ), .B(\un1_next_sum_iv_2[7] ), .C(sum_7), 
        .Y(N493));
    NOR2 inf_abs2_a_0_I_47 (.A(integral[21]), .B(integral[22]), .Y(
        \DWACT_FINC_E[11] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I89_Y (.A(N511), .B(N514), .Y(
        N639));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I10_P0N (.A(
        \un1_next_sum_iv_1[10] ), .B(\un1_next_sum_iv_2[10] ), .C(
        sum_10), .Y(N502));
    NOR2 inf_abs1_a_2_I_21 (.A(sr_new[6]), .B(sr_new[7]), .Y(
        \DWACT_FINC_E_0[3] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I5_G0N (.A(\i_adj[5]_net_1 ), 
        .B(\i_adj[7]_net_1 ), .Y(N281));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I176_Y (.A(\i_adj[18]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .C(N498), .Y(\next_ireg_3[22] ));
    NOR3 inf_abs2_a_0_I_8 (.A(integral[7]), .B(integral[6]), .C(
        integral[8]), .Y(N_24));
    XA1B \sumreg_RNO[16]  (.A(N1082), .B(ADD_40x40_fast_I434_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[16] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I383_Y_2 (.A(
        ADD_40x40_fast_I383_un1_Y_0), .B(N848), .C(
        ADD_40x40_fast_I383_Y_1), .Y(ADD_40x40_fast_I383_Y_2));
    NOR3B inf_abs2_a_0_I_19 (.A(\DWACT_FINC_E[2] ), .B(
        \DWACT_FINC_E_0[0] ), .C(integral[12]), .Y(N_20));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I78_Y (.A(I78_un1_Y), .B(N528_0), 
        .Y(N628));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I132_un1_Y (.A(N423), .B(N359), 
        .Y(I132_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I0_CO1 (.A(\i_adj[0]_net_1 ), 
        .B(\i_adj[2]_net_1 ), .Y(N266));
    OR2A un1_sumreg_0_0_ADD_40x40_fast_I26_P0N (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[26]_net_1 ), .Y(N550));
    NOR3B \ireg_RNI2LJQ[18]  (.A(\state[3]_net_1 ), .B(
        \ireg[18]_net_1 ), .C(integral_1_0), .Y(\ireg_m[18] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I229_Y (.A(N706), .B(N714), .Y(
        N788));
    XA1B \sumreg_RNO[13]  (.A(N1091), .B(ADD_40x40_fast_I431_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[13] ));
    XNOR2 inf_abs2_a_0_I_7 (.A(integral[8]), .B(N_25), .Y(
        \inf_abs2_a_0[2] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I133_un1_Y (.A(N425), .B(N266), 
        .Y(I133_un1_Y));
    XNOR2 inf_abs2_a_0_I_35 (.A(integral[18]), .B(N_15), .Y(
        \inf_abs2_a_0[12] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I1_P0N (.A(\i_adj[1]_net_1 ), .B(
        \i_adj[3]_net_1 ), .Y(N270));
    XOR2 inf_abs2_a_0_I_5 (.A(integral[6]), .B(integral[7]), .Y(
        \inf_abs2_a_0[1] ));
    OR2 \ireg_RNI6MRC2[25]  (.A(\un1_next_sum_0_iv_1[25] ), .B(
        \ireg_m[25] ), .Y(\un1_next_sum_0_iv[25] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I332_un1_Y (.A(N840), .B(N871), 
        .Y(I332_un1_Y));
    AND3 inf_abs2_a_0_I_61 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[15] ), .Y(N_6));
    AND3 inf_abs2_a_0_I_58 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[14] ), .Y(N_7));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I111_Y (.A(sum_2_d0), .B(sum_3), 
        .C(\un1_next_sum[0] ), .Y(N661));
    XA1B \sumreg_RNO[19]  (.A(N1073), .B(ADD_40x40_fast_I437_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[19] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I68_Y (.A(N341), .B(N338), .C(
        N337), .Y(N376));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I16_G0N (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(N519));
    XNOR2 inf_abs1_a_2_I_12 (.A(sr_new[4]), .B(N_10), .Y(
        \inf_abs1_a_2[4] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I446_Y_0 (.A(
        \sumreg[28]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I446_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I109_Y (.A(N391), .B(N383), .Y(
        N423));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I93_Y (.A(N505), .B(N508), .Y(
        N643));
    DFN1E1C0 \p_adj[12]  (.D(\inf_abs1_5[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[12]_net_1 ));
    DFN1E1C0 \p_adj[2]  (.D(\inf_abs1_5[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[2]_net_1 ));
    MX2 \i_adj_RNO[9]  (.A(integral[15]), .B(\inf_abs2_a_0[9] ), .S(
        integral[25]), .Y(\inf_abs2_5[9] ));
    DFN1E1C0 \ireg[18]  (.D(\next_ireg_3[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[18]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_1 (.A(N328), .B(N331), .C(
        ADD_22x22_fast_I143_Y_0), .Y(ADD_22x22_fast_I143_Y_1));
    NOR3A inf_abs2_a_0_I_13 (.A(\DWACT_FINC_E_0[0] ), .B(integral[9]), 
        .C(integral[10]), .Y(N_22));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I313_Y (.A(N816), .B(N800), .Y(
        N884));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I73_Y (.A(N538), .B(N535), .Y(
        N623));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_3 (.A(
        ADD_22x22_fast_I143_un1_Y_0), .B(N423), .C(
        ADD_22x22_fast_I143_Y_2), .Y(ADD_22x22_fast_I143_Y_3));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I45_Y (.A(\sumreg[35]_net_1 ), 
        .B(\sumreg[36]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N595)
        );
    DFN1E1C0 \ireg[9]  (.D(\next_ireg_3[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[9]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I382_Y_0 (.A(N679), .B(N687), .Y(
        ADD_40x40_fast_I382_Y_0));
    DFN1E1C0 \preg[14]  (.D(\p_adj[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[14]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I96_Y (.A(N498_0), .B(N502), .C(
        N501), .Y(N646));
    XNOR2 inf_abs2_a_0_I_59 (.A(integral[25]), .B(N_7), .Y(
        \inf_abs2_a_0[20] ));
    AND3 inf_abs2_a_0_I_24 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E_0[4] ));
    DFN1E1C0 \preg[9]  (.D(\p_adj[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[9]_net_1 ));
    AO1 \preg_RNI3S6D1[16]  (.A(\preg[16]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[16] ), .Y(
        \un1_next_sum_iv_1[16] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I426_Y_0 (.A(
        \un1_next_sum_iv_1[8] ), .B(\un1_next_sum_iv_2[8] ), .C(sum_8), 
        .Y(ADD_40x40_fast_I426_Y_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I379_Y (.A(I332_un1_Y), .B(
        ADD_40x40_fast_I379_Y_3), .C(I379_un1_Y), .Y(N1023));
    AO1 \preg_RNI707D1[18]  (.A(\preg[18]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[18] ), .Y(
        \un1_next_sum_iv_1[18] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I76_Y (.A(I76_un1_Y), .B(N531_0), 
        .Y(N626));
    DFN1P0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .PRE(n_rst_c), 
        .Q(sum_rdy));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I205_Y (.A(N690), .B(N682), .Y(
        N764));
    NOR2B inf_abs1_a_2_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_2));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I177_Y (.A(N653), .B(N649), .Y(
        N730));
    NOR3B inf_abs2_a_0_I_36 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .C(integral[18]), .Y(N_14));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I8_G0N (.A(
        \un1_next_sum_iv_1[8] ), .B(\un1_next_sum_iv_2[8] ), .C(sum_8), 
        .Y(N495));
    XA1B \sumreg_RNO[6]  (.A(N819), .B(ADD_40x40_fast_I424_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[6] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I218_un1_Y (.A(N703), .B(N696), 
        .Y(I218_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I71_Y (.A(N340), .B(N344), .Y(
        N379));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I350_Y_0 (.A(N793), .B(N778), .C(
        N777), .Y(ADD_40x40_fast_I350_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I145_Y (.A(N617), .B(N621), .Y(
        N698));
    AO1A \state_RNO[0]  (.A(sum_enable), .B(sum_rdy), .C(
        \state[5]_net_1 ), .Y(\state_ns[0] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I62_Y (.A(\sumreg[26]_net_1 ), 
        .B(\sumreg[27]_net_1 ), .C(\un1_next_sum_1_iv[26] ), .Y(N612));
    AO1 \preg_RNI1Q6D1[15]  (.A(\preg[15]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[15] ), .Y(
        \un1_next_sum_iv_1[15] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I380_Y (.A(N842), .B(N873), .C(
        ADD_40x40_fast_I380_Y_3), .Y(N1025));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I235_Y (.A(N712), .B(N720), .Y(
        N794));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I191_Y (.A(I116_un1_Y), .B(N664), 
        .Y(N745));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I455_Y_0 (.A(
        \sumreg[37]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I455_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I255_Y (.A(N740), .B(N732), .Y(
        N814));
    AO1 next_ireg_3_0_ADD_22x22_fast_I82_Y (.A(N355), .B(N352), .C(
        N351), .Y(N390));
    NOR2A inf_abs2_a_0_I_25 (.A(\DWACT_FINC_E_0[4] ), .B(integral[14]), 
        .Y(N_18));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I183_Y (.A(N659), .B(N655), .Y(
        N736));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I254_un1_Y (.A(N739), .B(N732), 
        .Y(I254_un1_Y));
    NOR3B \ireg_RNIHQKO[8]  (.A(integral_1_0), .B(\state[3]_net_1 ), 
        .C(\ireg[8]_net_1 ), .Y(\un3_next_sum_m[8] ));
    AO1 \preg_RNIPH6D1[11]  (.A(\preg[11]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[11] ), .Y(
        \un1_next_sum_iv_1[11] ));
    DFN1E1C0 \ireg[8]  (.D(\next_ireg_3[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[8]_net_1 ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I360_un1_Y (.A(N798), .B(N814), 
        .C(N666), .Y(I360_un1_Y));
    OA1 next_ireg_3_0_ADD_22x22_fast_I25_Y (.A(\i_adj[17]_net_1 ), .B(
        \i_adj[15]_net_1 ), .C(N315), .Y(N330));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I43_Y (.A(N285), .B(N288), .Y(
        N348));
    XNOR2 inf_abs1_a_2_I_35 (.A(sr_new[12]), .B(N_2), .Y(
        \inf_abs1_a_2[12] ));
    DFN1E1C0 \preg[8]  (.D(\p_adj[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[8]_net_1 ));
    XNOR2 inf_abs2_a_0_I_53 (.A(integral[24]), .B(N_9_0), .Y(
        \inf_abs2_a_0[18] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I301_Y (.A(N804), .B(N788), .Y(
        N872));
    DFN1E1C0 \i_adj[14]  (.D(\inf_abs2_5[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[14]_net_1 ));
    DFN1E1C0 \sumreg[32]  (.D(\next_sum[32] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(\sumreg[32]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I346_Y (.A(
        ADD_40x40_fast_I346_un1_Y_0), .B(N1085), .C(
        ADD_40x40_fast_I346_Y_0), .Y(N1037));
    AO1 next_ireg_3_0_ADD_22x22_fast_I28_Y (.A(N305), .B(N309), .C(
        N308), .Y(N333));
    NOR2A un1_sumreg_0_0_ADD_40x40_fast_I25_G0N (.A(\sumreg[25]_net_1 )
        , .B(\un1_next_sum_0_iv[25] ), .Y(N546));
    NOR3B \preg_RNIFEHP[12]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[12]_net_1 ), .Y(\un24_next_sum_m[12] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I249_Y (.A(N734), .B(N726), .Y(
        N808));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I351_Y (.A(
        ADD_40x40_fast_I351_un1_Y_0), .B(N1100), .C(
        ADD_40x40_fast_I351_Y_0), .Y(N1052));
    MX2 \i_adj_RNO[6]  (.A(integral[12]), .B(\inf_abs2_a_0[6] ), .S(
        integral[25]), .Y(\inf_abs2_5[6] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I188_Y (.A(N664), .B(N661), .C(
        N660), .Y(N741));
    AND3 inf_abs1_a_2_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(N_6_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I17_P0N (.A(
        \un1_next_sum_iv_1[17] ), .B(\un1_next_sum_iv_2[17] ), .C(
        sum_17), .Y(N523));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I16_P0N (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(N520));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I156_un1_Y (.A(N632), .B(N629), 
        .Y(I156_un1_Y));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I49_Y (.A(\sumreg[34]_net_1 ), 
        .B(\sumreg[33]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N599)
        );
    XNOR2 inf_abs2_a_0_I_26 (.A(integral[15]), .B(N_18), .Y(
        \inf_abs2_a_0[9] ));
    XA1B \sumreg_RNO[12]  (.A(N1094), .B(ADD_40x40_fast_I430_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[12] ));
    NOR2B \state_RNIL5TC[3]  (.A(\state[3]_net_1 ), .B(integral[25]), 
        .Y(next_sum_0_sqmuxa));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I54_Y (.A(\sumreg[30]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N604)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I315_Y (.A(N804), .B(N819), .C(
        N803), .Y(N1088));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I112_Y (.A(sum_1_d0), .B(
        sum_2_d0), .C(\un1_next_sum[0] ), .Y(N662));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I177_Y_0 (.A(\i_adj[19]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(ADD_22x22_fast_I177_Y_0));
    AO1 \preg_RNI5U6D1[17]  (.A(next_sum_1_sqmuxa_2), .B(
        \preg[17]_net_1 ), .C(\ireg_m[17] ), .Y(
        \un1_next_sum_iv_1[17] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I106_Y (.A(I106_un1_Y_0), .B(
        N486), .Y(N656));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I7_G0N (.A(
        \un1_next_sum_iv_1[7] ), .B(\un1_next_sum_iv_2[7] ), .C(sum_7), 
        .Y(N492_0));
    XA1 \ireg_RNIB94J[22]  (.A(integral_0_0), .B(\ireg[22]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[22] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I242_un1_Y (.A(N727), .B(N720), 
        .Y(I242_un1_Y));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I164_Y (.A(\i_adj[4]_net_1 ), .B(
        \i_adj[6]_net_1 ), .C(N394), .Y(\next_ireg_3[10] ));
    AO1 \preg_RNIVN6D1[14]  (.A(\preg[14]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[14] ), .Y(
        \un1_next_sum_iv_1[14] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_1 (.A(
        ADD_22x22_fast_I142_Y_0_a3_0), .B(N329), .C(
        ADD_22x22_fast_I142_Y_0_0), .Y(ADD_22x22_fast_I142_Y_0_1));
    XNOR2 inf_abs2_a_0_I_62 (.A(integral[25]), .B(N_6), .Y(
        \inf_abs2_a_0[21] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I419_Y_0 (.A(sum_1_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I419_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I68_Y (.A(N540), .B(N544), .C(
        N543), .Y(N618));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I22_G0N (.A(sum_22), .B(
        \un1_next_sum[22] ), .Y(N537));
    NOR2 inf_abs2_a_0_I_38 (.A(integral[18]), .B(integral[19]), .Y(
        \DWACT_FINC_E[8] ));
    NOR3 inf_abs2_a_0_I_41 (.A(integral[19]), .B(integral[18]), .C(
        integral[20]), .Y(\DWACT_FINC_E[9] ));
    MX2 \p_adj_RNO[9]  (.A(sr_new[9]), .B(\inf_abs1_a_2[9] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[9] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I136_Y (.A(N612), .B(N608), .Y(
        N689));
    DFN1E1C0 \sumreg[33]  (.D(\next_sum[33] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(\sumreg[33]_net_1 ));
    XA1B \sumreg_RNO[2]  (.A(N745), .B(ADD_40x40_fast_I420_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[2] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I156_Y (.A(I156_un1_Y), .B(N628), 
        .Y(N709));
    NOR3B \ireg_RNITG4H[6]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[6]_net_1 ), .C(integral_0_0), .Y(\ireg_m[6] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I352_un1_Y_0 (.A(N798), .B(
        N782), .Y(ADD_40x40_fast_I352_un1_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I100_Y (.A(N492_0), .B(N496), .C(
        N495), .Y(N650));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I165_Y_0 (.A(\i_adj[7]_net_1 ), 
        .B(\i_adj[5]_net_1 ), .Y(ADD_22x22_fast_I165_Y_0));
    DFN1E1C0 \i_adj[12]  (.D(\inf_abs2_5[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[12]_net_1 ));
    NOR2B \i_adj_RNO[19]  (.A(\inf_abs2_a_0[19] ), .B(integral[25]), 
        .Y(\inf_abs2_5[19] ));
    NOR3B \ireg_RNIVEDM[16]  (.A(integral_0_0), .B(\state[3]_net_1 ), 
        .C(\ireg[16]_net_1 ), .Y(\un3_next_sum_m[16] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I359_un1_Y (.A(N796), .B(N812), 
        .C(N745), .Y(I359_un1_Y));
    OA1 next_ireg_3_0_ADD_22x22_fast_I39_Y (.A(\i_adj[8]_net_1 ), .B(
        \i_adj[10]_net_1 ), .C(N294), .Y(N344));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I143_un1_Y_0 (.A(N375), .B(N367)
        , .C(N359), .Y(ADD_22x22_fast_I143_un1_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y_0 (.A(N335), .B(N332), .C(
        N331), .Y(ADD_22x22_fast_I126_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I14_G0N (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .Y(N308));
    DFN1E1C0 \sumreg[30]  (.D(\next_sum[30] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(\sumreg[30]_net_1 ));
    AND3 inf_abs2_a_0_I_39 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E_0[7] ), .C(\DWACT_FINC_E[8] ), .Y(N_13));
    AO1 next_ireg_3_0_ADD_22x22_fast_I24_Y (.A(N311), .B(N315), .C(
        N314), .Y(N329));
    OA1 next_ireg_3_0_ADD_22x22_fast_I37_Y (.A(\i_adj[12]_net_1 ), .B(
        \i_adj[10]_net_1 ), .C(N294), .Y(N342));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I302_Y (.A(N805), .B(N790), .C(
        N789), .Y(N873));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I292_un1_Y (.A(N706), .B(N698), 
        .C(N795), .Y(I292_un1_Y));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I130_Y (.A(N606), .B(N602), .Y(
        N683));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I80_Y (.A(N522_0), .B(N526), .C(
        N525_0), .Y(N630));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I346_un1_Y_0 (.A(N786), .B(
        N770), .Y(ADD_40x40_fast_I346_un1_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I0_G0N (.A(N_228), .B(sum_0_d0)
        , .Y(N471));
    NOR3B \ireg_RNI1KJQ[17]  (.A(\state[3]_net_1 ), .B(
        \ireg[17]_net_1 ), .C(integral_1_0), .Y(\ireg_m[17] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I150_Y (.A(I150_un1_Y), .B(N622), 
        .Y(N703));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I161_Y (.A(N633), .B(N637), .Y(
        N714));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I40_Y (.A(N287), .B(
        \i_adj[8]_net_1 ), .C(\i_adj[10]_net_1 ), .Y(N345));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I172_Y_0 (.A(\i_adj[12]_net_1 ), 
        .B(\i_adj[14]_net_1 ), .Y(ADD_22x22_fast_I172_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I346_Y_0 (.A(N785), .B(N770), .C(
        N769), .Y(ADD_40x40_fast_I346_Y_0));
    OR3 \preg_RNIPKEQ1[17]  (.A(\un24_next_sum_m[17] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[17] ), .Y(
        \un1_next_sum_iv_2[17] ));
    OA1A un1_sumreg_0_0_ADD_40x40_fast_I63_Y (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[27]_net_1 ), .C(N550), .Y(
        N613));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I187_Y (.A(
        ADD_40x40_fast_I187_Y_0), .B(N659), .Y(N740));
    XA1B \sumreg_RNO[4]  (.A(N823), .B(ADD_40x40_fast_I422_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[4] ));
    NOR3B \preg_RNIGFHP[13]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[13]_net_1 ), .Y(\un24_next_sum_m[13] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I352_Y (.A(I294_un1_Y), .B(N781), 
        .C(I352_un1_Y), .Y(N1055));
    XA1B \sumreg_RNO[5]  (.A(N821), .B(ADD_40x40_fast_I423_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[5] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I378_Y (.A(
        ADD_40x40_fast_I378_Y_3), .B(I378_un1_Y), .C(I330_un1_Y), .Y(
        N1021));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I45_Y (.A(N282), .B(N285), .Y(
        N350));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I171_Y (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .C(N513), .Y(\next_ireg_3[17] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_o3_0_0 (.A(N337), .B(
        N334), .C(N333), .Y(ADD_22x22_fast_I142_Y_0_o3_0_0));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I432_Y_0 (.A(
        \un1_next_sum_iv_1[14] ), .B(\un1_next_sum_iv_2[14] ), .C(
        sum_14), .Y(ADD_40x40_fast_I432_Y_0));
    DFN1E1C0 \sumreg[37]  (.D(\next_sum[37] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(\sumreg[37]_net_1 ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I51_Y (.A(\sumreg[33]_net_1 ), 
        .B(\sumreg[32]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N601)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I383_Y_1 (.A(N764), .B(N779), .C(
        ADD_40x40_fast_I383_Y_0), .Y(ADD_40x40_fast_I383_Y_1));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I23_P0N (.A(\un1_next_sum[23] ), 
        .B(sum_23), .Y(N541));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_2 (.A(N367), .B(N374), .C(
        ADD_22x22_fast_I143_Y_1), .Y(ADD_22x22_fast_I143_Y_2));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I66_Y (.A(N543), .B(N547), .C(
        N546), .Y(N616));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I445_Y_0 (.A(
        \sumreg[27]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I445_Y_0));
    NOR3B \ireg_RNI963J[11]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[11]_net_1 ), .Y(\un3_next_sum_m[11] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I109_Y (.A(N481), .B(N484), .Y(
        N659));
    XNOR2 inf_abs2_a_0_I_28 (.A(integral[16]), .B(N_17), .Y(
        \inf_abs2_a_0[10] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I19_P0N (.A(\un1_next_sum[19] ), 
        .B(sum_19), .Y(N529));
    NOR3 inf_abs2_a_0_I_33 (.A(integral[16]), .B(integral[15]), .C(
        integral[17]), .Y(\DWACT_FINC_E_0[7] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I55_Y (.A(\sumreg[30]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N605)
        );
    DFN1C0 \state_1[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_1[2]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I48_Y (.A(N275), .B(N279), .C(
        N278), .Y(N353));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I3_G0N (.A(sum_3), .B(
        \un1_next_sum[0] ), .Y(N480));
    MX2 \i_adj_RNO[4]  (.A(integral[10]), .B(\inf_abs2_a_0[4] ), .S(
        integral[25]), .Y(\inf_abs2_5[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I210_Y (.A(N695), .B(N688), .C(
        N687), .Y(N769));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I15_G0N (.A(
        \un1_next_sum_iv_1[15] ), .B(\un1_next_sum_iv_2[15] ), .C(
        sum_15), .Y(N516));
    NOR3B \ireg_RNIC93J[14]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[14]_net_1 ), .Y(\un3_next_sum_m[14] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I425_Y_0 (.A(
        \un1_next_sum_iv_1[7] ), .B(\un1_next_sum_iv_2[7] ), .C(sum_7), 
        .Y(ADD_40x40_fast_I425_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I139_Y (.A(N611), .B(N615), .Y(
        N692));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I277_Y (.A(N706), .B(N698), .C(
        N764), .Y(N848));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I159_Y (.A(N635), .B(N631), .Y(
        N712));
    DFN1E1C0 \i_adj[13]  (.D(\inf_abs2_5[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[13]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I104_Y (.A(N486), .B(N490), .C(
        N489), .Y(N654));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I115_un1_Y (.A(N393), .B(N266), 
        .Y(I115_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I54_un1_Y (.A(N270), .B(N266), 
        .Y(I54_un1_Y));
    NOR3 inf_abs2_a_0_I_29 (.A(integral[12]), .B(integral[14]), .C(
        integral[13]), .Y(\DWACT_FINC_E[5] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I130_Y_0 (.A(N386), .B(N379), .C(
        N378), .Y(ADD_22x22_fast_I130_Y_0));
    DFN1E1C0 \preg[12]  (.D(\p_adj[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[12]_net_1 ));
    MX2 \i_adj_RNO[2]  (.A(integral[8]), .B(\inf_abs2_a_0[2] ), .S(
        integral[25]), .Y(\inf_abs2_5[2] ));
    DFN1E1C0 \i_adj[5]  (.D(\inf_abs2_5[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[5]_net_1 ));
    DFN1E1C0 \ireg[20]  (.D(\next_ireg_3[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[20]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I379_Y_0 (.A(\sumreg[36]_net_1 )
        , .B(\sumreg[37]_net_1 ), .C(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I379_Y_0));
    OR3 un1_sumreg_0_0_ADD_m8_i_o4_1 (.A(sum_2_d0), .B(sum_1_d0), .C(
        sum_0_d0), .Y(ADD_m8_i_o4_1));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I378_Y_0 (.A(\sumreg[38]_net_1 )
        , .B(\sumreg[37]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(
        ADD_40x40_fast_I378_Y_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I380_Y_3 (.A(I270_un1_Y), .B(
        ADD_40x40_fast_I380_Y_1), .C(I380_un1_Y), .Y(
        ADD_40x40_fast_I380_Y_3));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I134_Y (.A(N610), .B(N606), .Y(
        N687));
    DFN1E1C0 \i_adj[0]  (.D(\inf_abs2_5[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[0]_net_1 ));
    DFN1E1C0 \p_adj[6]  (.D(\inf_abs1_5[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[6]_net_1 ));
    MX2 \p_adj_RNO[4]  (.A(sr_new[4]), .B(\inf_abs1_a_2[4] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I154_Y (.A(N630), .B(N627), .C(
        N626), .Y(N707));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I211_Y (.A(N688), .B(N696), .Y(
        N770));
    XA1 \ireg_RNIA84J[21]  (.A(integral_0_0), .B(\ireg[21]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[21] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I270_un1_Y (.A(N758), .B(N773), 
        .Y(I270_un1_Y));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I12_G0N (.A(
        \un1_next_sum_iv_1[12] ), .B(\un1_next_sum_iv_2[12] ), .C(
        sum_12), .Y(N507_0));
    XA1B \sumreg_RNO[24]  (.A(N1058), .B(ADD_40x40_fast_I442_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[24] ));
    NOR3B \ireg_RNI853J[10]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[10]_net_1 ), .Y(\un3_next_sum_m[10] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I59_Y (.A(N328), .B(N332), .Y(
        N367));
    MX2 \i_adj_RNO[0]  (.A(integral[6]), .B(integral[6]), .S(
        integral[25]), .Y(\inf_abs2_5[0] ));
    OR3 \ireg_RNIIJ171[23]  (.A(next_sum_0_sqmuxa_2), .B(
        next_sum_0_sqmuxa_1), .C(\un1_next_sum_iv_0[23] ), .Y(
        \un1_next_sum[23] ));
    AND3 inf_abs2_a_0_I_42 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E_0[7] ), .C(\DWACT_FINC_E[9] ), .Y(N_12_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I17_P0N_i_o3 (.A(
        \i_adj[19]_net_1 ), .B(\i_adj[17]_net_1 ), .Y(N_9));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I218_Y (.A(I218_un1_Y), .B(N695), 
        .Y(N777));
    XNOR2 inf_abs2_a_0_I_23 (.A(integral[14]), .B(N_19), .Y(
        \inf_abs2_a_0[8] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I66_Y (.A(N339), .B(N336), .C(
        N335), .Y(N374));
    AO1 \preg_RNILUE71[9]  (.A(\preg[9]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[9] ), .Y(
        \un1_next_sum_iv_1[9] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I44_Y (.A(N281), .B(N285), .C(
        N284), .Y(N349));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I439_Y_0 (.A(sum_21), .B(
        \un1_next_sum[21] ), .Y(ADD_40x40_fast_I439_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I450_Y_0 (.A(
        \sumreg[32]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I450_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I234_Y (.A(N719), .B(N712), .C(
        N711), .Y(N793));
    NOR3 inf_abs1_a_2_I_33 (.A(sr_new[10]), .B(sr_new[9]), .C(
        sr_new[11]), .Y(\DWACT_FINC_E[7] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I384_Y (.A(N850), .B(N881), .C(
        ADD_40x40_fast_I384_Y_2), .Y(N1033));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I254_Y (.A(I254_un1_Y), .B(N731), 
        .Y(N813));
    MX2 \i_adj_RNO[7]  (.A(integral[13]), .B(\inf_abs2_a_0[7] ), .S(
        integral[25]), .Y(\inf_abs2_5[7] ));
    DFN1E1C0 \i_adj[21]  (.D(\inf_abs2_5[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[21]_net_1 ));
    XA1B \sumreg_RNO[9]  (.A(N1103), .B(ADD_40x40_fast_I427_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[9] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I59_Y (.A(\sumreg[29]_net_1 ), 
        .B(\sumreg[28]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N609)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I162_Y (.A(N638), .B(N635), .C(
        N634), .Y(N715));
    NOR3A \state_RNI9POH[4]  (.A(integral_1_0), .B(\state[5]_net_1 ), 
        .C(\state[4]_net_1 ), .Y(N_232));
    NOR2A \state_RNIL5TC_0[3]  (.A(\state[3]_net_1 ), .B(integral[25]), 
        .Y(next_sum_1_sqmuxa));
    DFN1E1C0 \ireg[14]  (.D(\next_ireg_3[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[14]_net_1 ));
    DFN1E1C0 \p_adj[11]  (.D(\inf_abs1_5[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[11]_net_1 ));
    OR3 \ireg_RNIMFCG1[25]  (.A(next_sum_1_sqmuxa_2), .B(
        next_sum_1_sqmuxa_1), .C(\un3_next_sum_m[25] ), .Y(
        \un1_next_sum_0_iv_1[25] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I82_Y (.A(N519), .B(N523), .C(
        N522_0), .Y(N632));
    DFN1E1C0 \i_adj[16]  (.D(\inf_abs2_5[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[16]_net_1 ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I4_P0N (.A(\i_adj[4]_net_1 ), .B(
        \i_adj[6]_net_1 ), .Y(N279));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I178_Y_0 (.A(\i_adj[20]_net_1 ), 
        .B(\i_adj[18]_net_1 ), .Y(ADD_22x22_fast_I178_Y_0));
    NOR3B \ireg_RNIRDJQ[11]  (.A(\state[3]_net_1 ), .B(
        \ireg[11]_net_1 ), .C(integral_1_0), .Y(\ireg_m[11] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I131_Y_0 (.A(N345), .B(N342), .C(
        N341), .Y(ADD_22x22_fast_I131_Y_0));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I437_Y_0 (.A(sum_19), .B(
        \un1_next_sum[19] ), .Y(ADD_40x40_fast_I437_Y_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I13_P0N (.A(
        \un1_next_sum_iv_1[13] ), .B(\un1_next_sum_iv_2[13] ), .C(
        sum_13), .Y(N511));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I32_Y (.A(N299), .B(
        \i_adj[12]_net_1 ), .C(\i_adj[14]_net_1 ), .Y(N337));
    MX2 \i_adj_RNO[11]  (.A(integral[17]), .B(\inf_abs2_a_0[11] ), .S(
        integral_1_0), .Y(\inf_abs2_5[11] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I15_G0N (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(N311));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I385_Y_2 (.A(I280_un1_Y), .B(
        ADD_40x40_fast_I385_Y_0), .C(I385_un1_Y), .Y(
        ADD_40x40_fast_I385_Y_2));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I298_Y (.A(N801), .B(N786), .C(
        N785), .Y(N869));
    DFN1E1C0 \ireg[4]  (.D(\i_adj[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[4]_net_1 ));
    OR2 \preg_RNI4FL33[6]  (.A(\un1_next_sum_iv_2[6] ), .B(
        \un1_next_sum_iv_1[6] ), .Y(\un1_next_sum[6] ));
    MX2 \p_adj_RNO[11]  (.A(sr_new[11]), .B(\inf_abs1_a_2[11] ), .S(
        sr_new_1_0), .Y(\inf_abs1_5[11] ));
    AX1D next_ireg_3_0_ADD_22x22_fast_I172_Y (.A(I130_un1_Y), .B(
        ADD_22x22_fast_I130_Y_0), .C(ADD_22x22_fast_I172_Y_0), .Y(
        \next_ireg_3[18] ));
    XA1B \sumreg_RNO[37]  (.A(N1025), .B(ADD_40x40_fast_I455_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[37] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I381_un1_Y (.A(N876), .B(N823), 
        .C(N844), .Y(I381_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I141_Y (.A(N613), .B(N617), .Y(
        N694));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I83_Y (.A(N356), .B(N352), .Y(
        N391));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I111_Y (.A(N393), .B(N385), .Y(
        N425));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I175_Y (.A(N651), .B(N647), .Y(
        N728));
    AO1 \preg_RNIHQE71[7]  (.A(\preg[7]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[7] ), .Y(
        \un1_next_sum_iv_1[7] ));
    NOR3B \ireg_RNIFOKO[6]  (.A(integral_1_0), .B(\state[3]_net_1 ), 
        .C(\ireg[6]_net_1 ), .Y(\un3_next_sum_m[6] ));
    DFN1E1C0 \sumreg[24]  (.D(\next_sum[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[24]_net_1 ));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I26_Y (.A(N308), .B(
        \i_adj[17]_net_1 ), .C(\i_adj[15]_net_1 ), .Y(N331));
    XA1 \ireg_RNICA4J[23]  (.A(integral_0_0), .B(\ireg[23]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[23] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I24_G0N (.A(\un1_next_sum[24] )
        , .B(\sumreg[24]_net_1 ), .Y(N543));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I175_Y (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .C(N_11), .Y(\next_ireg_3[21] ));
    NOR3 \state_RNIG3OG[6]  (.A(sum_rdy), .B(\state[6]_net_1 ), .C(
        \state_0[1]_net_1 ), .Y(N_416_0));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I431_Y_0 (.A(
        \un1_next_sum_iv_1[13] ), .B(\un1_next_sum_iv_2[13] ), .C(
        sum_13), .Y(ADD_40x40_fast_I431_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I300_Y (.A(N803), .B(N788), .C(
        N787), .Y(N871));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I103_Y (.A(N490), .B(N493), .Y(
        N653));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I88_Y (.A(N510), .B(N514), .C(
        N513_0), .Y(N638));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I0_P0N (.A(N_228), .B(sum_0_d0), 
        .Y(N472));
    NOR2B \state_RNI1OD9[5]  (.A(\state[5]_net_1 ), .B(sr_new[12]), .Y(
        next_sum_0_sqmuxa_2));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I260_Y (.A(N740), .B(N666), .C(
        N739), .Y(N821));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I8_P0N (.A(
        \un1_next_sum_iv_1[8] ), .B(\un1_next_sum_iv_2[8] ), .C(sum_8), 
        .Y(N496));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I106_un1_Y (.A(N483), .B(N487), 
        .Y(I106_un1_Y_0));
    MX2 \i_adj_RNO[15]  (.A(integral[21]), .B(\inf_abs2_a_0[15] ), .S(
        integral_1_0), .Y(\inf_abs2_5[15] ));
    DFN1E1C0 \sumreg[14]  (.D(\next_sum[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_14));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I350_Y (.A(
        ADD_40x40_fast_I350_un1_Y_0), .B(N1097), .C(
        ADD_40x40_fast_I350_Y_0), .Y(N1049));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I203_Y (.A(N680), .B(N688), .Y(
        N762));
    NOR2B \i_adj_RNO[20]  (.A(\inf_abs2_a_0[20] ), .B(integral[25]), 
        .Y(\inf_abs2_5[20] ));
    XNOR2 inf_abs1_a_2_I_14 (.A(sr_new[5]), .B(N_9_1), .Y(
        \inf_abs1_a_2[5] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I170_Y_0 (.A(\i_adj[12]_net_1 ), 
        .B(\i_adj[10]_net_1 ), .Y(ADD_22x22_fast_I170_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I133_Y (.A(N609), .B(N605), .Y(
        N686));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I215_Y (.A(N700), .B(N692), .Y(
        N774));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I279_Y (.A(N766), .B(N782), .Y(
        N850));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I153_Y (.A(N625), .B(N629), .Y(
        N706));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I79_Y (.A(N352), .B(N348), .Y(
        N387));
    XA1B \sumreg_RNO[30]  (.A(N1040), .B(ADD_40x40_fast_I448_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[30] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I77_Y (.A(N350), .B(N346), .Y(
        N385));
    NOR2B \state_RNI5HFA[4]  (.A(derivative_0), .B(\state[4]_net_1 ), 
        .Y(next_sum_0_sqmuxa_1));
    XNOR2 inf_abs2_a_0_I_9 (.A(integral[9]), .B(N_24), .Y(
        \inf_abs2_a_0[3] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I233_Y (.A(N710), .B(N718), .Y(
        N792));
    XA1B \sumreg_RNO[31]  (.A(N1037), .B(ADD_40x40_fast_I449_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[31] ));
    NOR3 inf_abs2_a_0_I_10 (.A(integral[7]), .B(integral[6]), .C(
        integral[8]), .Y(\DWACT_FINC_E_0[0] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I440_Y_0 (.A(sum_22), .B(
        \un1_next_sum[22] ), .Y(ADD_40x40_fast_I440_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I253_Y (.A(N738), .B(N730), .Y(
        N812));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I52_Y (.A(N269), .B(
        \i_adj[2]_net_1 ), .C(\i_adj[4]_net_1 ), .Y(N357));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I108_Y (.A(N480), .B(N484), .C(
        N483), .Y(N658));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I261_Y (.A(I116_un1_Y), .B(N741), 
        .Y(N823));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I173_Y (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[15]_net_1 ), .C(N507), .Y(\next_ireg_3[19] ));
    OR3 \ireg_RNIHI171[22]  (.A(next_sum_0_sqmuxa_2), .B(
        next_sum_0_sqmuxa_1), .C(\un1_next_sum_iv_0[22] ), .Y(
        \un1_next_sum[22] ));
    NOR2 inf_abs1_a_2_I_15 (.A(sr_new[4]), .B(sr_new[3]), .Y(
        \DWACT_FINC_E_0[1] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I83_Y (.A(N523), .B(N520), .Y(
        N633));
    XA1B \sumreg_RNO[25]  (.A(N1055), .B(ADD_40x40_fast_I443_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[25] ));
    DFN1E1C0 \i_adj[11]  (.D(\inf_abs2_5[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[11]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I307_Y (.A(N810), .B(N794), .Y(
        N878));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I138_Y (.A(N614), .B(N611), .C(
        N610), .Y(N691));
    DFN1E1C0 \ireg[11]  (.D(\next_ireg_3[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[11]_net_1 ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I420_Y_0 (.A(sum_2_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I420_Y_0));
    DFN1C0 \state[3]  (.D(\state[6]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[3]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I158_Y (.A(N634), .B(N631), .C(
        N630), .Y(N711));
    NOR3B \ireg_RNIIRKO[9]  (.A(integral_1_0), .B(\state[3]_net_1 ), 
        .C(\ireg[9]_net_1 ), .Y(\un3_next_sum_m[9] ));
    MX2 \i_adj_RNO[17]  (.A(integral[23]), .B(\inf_abs2_a_0[17] ), .S(
        integral_1_0), .Y(\inf_abs2_5[17] ));
    DFN1E1C0 \i_adj[1]  (.D(\inf_abs2_5[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[1]_net_1 ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I80_Y (.A(I80_un1_Y), .B(N349), 
        .Y(N388));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I86_Y (.A(N513_0), .B(N517), .C(
        N516), .Y(N636));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I236_Y (.A(N721), .B(N714), .C(
        N713), .Y(N795));
    DFN1E1C0 \sumreg[3]  (.D(\next_sum[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNI172K[6]_net_1 ), .Q(sum_3));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I220_Y (.A(N705), .B(N698), .C(
        N697), .Y(N779));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I256_Y (.A(N741), .B(N734), .C(
        N733), .Y(N815));
    DFN1E1C0 \sumreg_1[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(sum_1_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I4_G0N (.A(\i_adj[4]_net_1 ), 
        .B(\i_adj[6]_net_1 ), .Y(N278));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I357_Y (.A(N876), .B(N823), .C(
        N875), .Y(N1070));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I85_Y (.A(
        ADD_22x22_fast_I85_Y_0), .B(N354), .Y(N393));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I24_P0N (.A(\un1_next_sum[24] ), 
        .B(\sumreg[24]_net_1 ), .Y(N544));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I142_Y (.A(N618), .B(N615), .C(
        N614), .Y(N695));
    DFN1C0 \state_0[1]  (.D(\state_RNIK76G[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_0[1]_net_1 ));
    NOR3 inf_abs2_a_0_I_50 (.A(integral[22]), .B(integral[21]), .C(
        integral[23]), .Y(\DWACT_FINC_E[12] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I347_un1_Y_0 (.A(N788), .B(
        N772), .Y(ADD_40x40_fast_I347_un1_Y_0));
    AO1 \preg_RNIFOE71[6]  (.A(\preg[6]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[6] ), .Y(
        \un1_next_sum_iv_1[6] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I3_G0N (.A(\i_adj[3]_net_1 ), 
        .B(\i_adj[5]_net_1 ), .Y(N275));
    XNOR2 inf_abs1_a_2_I_9 (.A(sr_new[3]), .B(N_11_1), .Y(
        \inf_abs1_a_2[3] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I74_un1_Y (.A(N531_0), .B(N535)
        , .Y(I74_un1_Y));
    NOR3B inf_abs1_a_2_I_16 (.A(\DWACT_FINC_E_0[1] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[5]), .Y(N_8_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I46_Y (.A(N278), .B(N282), .C(
        N281), .Y(N351));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I13_G0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[15]_net_1 ), .Y(N305));
    VCC VCC_i (.Y(VCC));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I14_G0N (.A(
        \un1_next_sum_iv_1[14] ), .B(\un1_next_sum_iv_2[14] ), .C(
        sum_14), .Y(N513_0));
    AO1 \preg_RNIJSE71[8]  (.A(\preg[8]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[8] ), .Y(
        \un1_next_sum_iv_1[8] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I116_Y (.A(N471), .B(I116_un1_Y), 
        .Y(N666));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I50_Y (.A(\sumreg[32]_net_1 ), 
        .B(\sumreg[33]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N600)
        );
    AND3 inf_abs1_a_2_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(
        \DWACT_FINC_E[4] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I6_G0N (.A(\un1_next_sum[6] ), 
        .B(sum_6), .Y(N489));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I185_Y (.A(N661), .B(N657), .Y(
        N738));
    OA1 next_ireg_3_0_ADD_22x22_fast_I85_Y_0 (.A(\i_adj[2]_net_1 ), .B(
        \i_adj[4]_net_1 ), .C(N270), .Y(ADD_22x22_fast_I85_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I448_Y_0 (.A(
        \sumreg[30]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I448_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I107_Y (.A(N484), .B(N487), .Y(
        N657));
    AO1 next_ireg_3_0_ADD_22x22_fast_I129_Y_0 (.A(N384), .B(N377), .C(
        N376), .Y(ADD_22x22_fast_I129_Y_0));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I130_un1_Y (.A(N379), .B(N387), 
        .C(N394), .Y(I130_un1_Y));
    AO1 next_ireg_3_0_ADD_22x22_fast_I112_Y (.A(N387), .B(N394), .C(
        N386), .Y(N522));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I228_Y (.A(N713), .B(N706), .C(
        N705), .Y(N787));
    NOR3 inf_abs1_a_2_I_8 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2]), 
        .Y(N_11_1));
    XA1B \sumreg_RNO[26]  (.A(N1052), .B(ADD_40x40_fast_I444_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[26] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I454_Y_0 (.A(
        \sumreg[36]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I454_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I110_Y (.A(sum_2_d0), .B(
        \un1_next_sum[0] ), .C(N480), .Y(N660));
    XA1B \sumreg_RNO[17]  (.A(N1079), .B(ADD_40x40_fast_I435_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[17] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I359_Y (.A(N879), .B(I359_un1_Y), 
        .Y(N1076));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I137_Y (.A(N613), .B(N609), .Y(
        N690));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I129_un1_Y_0 (.A(N377), .B(N385)
        , .Y(ADD_22x22_fast_I129_un1_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I453_Y_0 (.A(
        \sumreg[35]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I453_Y_0));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I48_Y (.A(\sumreg[33]_net_1 ), 
        .B(\sumreg[34]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(
        I122_un1_Y));
    NOR2A inf_abs1_a_2_I_25 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .Y(
        N_5));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I157_Y (.A(N629), .B(N633), .Y(
        N710));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I428_Y_0 (.A(
        \un1_next_sum_iv_1[10] ), .B(\un1_next_sum_iv_2[10] ), .C(
        sum_10), .Y(ADD_40x40_fast_I428_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I312_Y (.A(N815), .B(N800), .C(
        N799), .Y(N883));
    DFN1E1C0 \preg[11]  (.D(\p_adj[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[11]_net_1 ));
    XA1B \sumreg_RNO[23]  (.A(N1061), .B(ADD_40x40_fast_I441_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[23] ));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I131_un1_Y (.A(N389), .B(N381), 
        .C(N396), .Y(I131_un1_Y));
    DFN1E1C0 \sumreg[22]  (.D(\next_sum[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_22));
    OR2 next_ireg_3_0_ADD_22x22_fast_I115_Y (.A(I115_un1_Y), .B(N392), 
        .Y(N531));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I5_P0N (.A(\un1_next_sum[5] ), 
        .B(sum_5), .Y(N487));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I20_G0N (.A(\un1_next_sum[20] )
        , .B(sum_20), .Y(N531_0));
    DFN1E1C0 \ireg[13]  (.D(\next_ireg_3[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[13]_net_1 ));
    XA1B \sumreg_RNO[29]  (.A(N1043), .B(ADD_40x40_fast_I447_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[29] ));
    DFN1E1C0 \p_adj[8]  (.D(\inf_abs1_5[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[8]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I61_Y (.A(N330), .B(N334), .Y(
        N369));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I351_Y_0 (.A(N779), .B(
        I292_un1_Y), .Y(ADD_40x40_fast_I351_Y_0));
    OR3 \ireg_RNIFG171[20]  (.A(next_sum_0_sqmuxa_2), .B(
        next_sum_0_sqmuxa_1), .C(\un1_next_sum_iv_0[20] ), .Y(
        \un1_next_sum[20] ));
    AX1D next_ireg_3_0_ADD_22x22_fast_I177_Y (.A(I124_un1_Y), .B(
        ADD_22x22_fast_I144_Y_2), .C(ADD_22x22_fast_I177_Y_0), .Y(
        \next_ireg_3[23] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I84_Y (.A(N357), .B(N354), .C(
        N353), .Y(N392));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I240_Y (.A(N725), .B(N718), .C(
        N717), .Y(N799));
    XNOR2 inf_abs1_a_2_I_7 (.A(sr_new[2]), .B(N_12), .Y(
        \inf_abs1_a_2[2] ));
    XNOR2 inf_abs2_a_0_I_17 (.A(integral[12]), .B(N_21), .Y(
        \inf_abs2_a_0[6] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_1_1 (.A(
        \i_adj[19]_net_1 ), .B(\i_adj[17]_net_1 ), .Y(N_14_1));
    DFN1E1C0 \sumreg[12]  (.D(\next_sum[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_12));
    DFN1E1C0 \ireg[15]  (.D(\next_ireg_3[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[15]_net_1 ));
    XA1B \sumreg_RNO[1]  (.A(N666), .B(ADD_40x40_fast_I419_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[1] ));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I179_Y (.A(\i_adj[19]_net_1 ), 
        .B(\i_adj[21]_net_1 ), .C(N492), .Y(\next_ireg_3[25] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I97_Y (.A(N502), .B(N499), .Y(
        N647));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I280_un1_Y (.A(N768), .B(N783), 
        .Y(I280_un1_Y));
    DFN1E1C0 \sumreg_2[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI172K[6]_net_1 ), .Q(sum_2_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I7_P0N (.A(\i_adj[7]_net_1 ), .B(
        \i_adj[9]_net_1 ), .Y(N288));
    NOR3 inf_abs1_a_2_I_18 (.A(sr_new[5]), .B(sr_new[4]), .C(sr_new[3])
        , .Y(\DWACT_FINC_E_0[2] ));
    XNOR2 inf_abs1_a_2_I_26 (.A(sr_new[9]), .B(N_5), .Y(
        \inf_abs1_a_2[9] ));
    
endmodule


module sig_gen_3(
       vd_done,
       n_rst_c,
       clk_c,
       vd_rdy
    );
input  vd_done;
input  n_rst_c;
input  clk_c;
output vd_rdy;

    wire sig_prev_i, sig_prev_net_1, sig_old_i_0, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(clk_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev (.D(vd_done), .CLK(clk_c), .CLR(n_rst_c), .Q(
        sig_prev_net_1));
    INV sig_old_RNO (.A(sig_prev_net_1), .Y(sig_prev_i));
    NOR2B sig_old_RNIO2D5 (.A(sig_prev_net_1), .B(sig_old_i_0), .Y(
        vd_rdy));
    GND GND_i (.Y(GND));
    
endmodule


module spi_stp_12s_1_6_0(
       cur_vd,
       N_29,
       din_fb_c,
       n_rst_c,
       sck_33_c
    );
output [11:0] cur_vd;
input  N_29;
input  din_fb_c;
input  n_rst_c;
input  sck_33_c;

    wire GND, VCC;
    
    DFN1E0C0 \sr[7]  (.D(cur_vd[6]), .CLK(sck_33_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[7]));
    DFN1E0C0 \sr[5]  (.D(cur_vd[4]), .CLK(sck_33_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[5]));
    DFN1E0C0 \sr[10]  (.D(cur_vd[9]), .CLK(sck_33_c), .CLR(n_rst_c), 
        .E(N_29), .Q(cur_vd[10]));
    DFN1E0C0 \sr[8]  (.D(cur_vd[7]), .CLK(sck_33_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[8]));
    DFN1E0C0 \sr[3]  (.D(cur_vd[2]), .CLK(sck_33_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[3]));
    DFN1E0C0 \sr[1]  (.D(cur_vd[0]), .CLK(sck_33_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[1]));
    DFN1E0C0 \sr[2]  (.D(cur_vd[1]), .CLK(sck_33_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[2]));
    DFN1E0C0 \sr[9]  (.D(cur_vd[8]), .CLK(sck_33_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[9]));
    VCC VCC_i (.Y(VCC));
    DFN1E0C0 \sr[11]  (.D(cur_vd[10]), .CLK(sck_33_c), .CLR(n_rst_c), 
        .E(N_29), .Q(cur_vd[11]));
    DFN1E0C0 \sr[0]  (.D(din_fb_c), .CLK(sck_33_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[0]));
    GND GND_i (.Y(GND));
    DFN1E0C0 \sr[6]  (.D(cur_vd[5]), .CLK(sck_33_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[6]));
    DFN1E0C0 \sr[4]  (.D(cur_vd[3]), .CLK(sck_33_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[4]));
    
endmodule


module sig_gen_0_0(
       cs_i_1,
       n_rst_c,
       sck_33_c,
       vd_done
    );
input  cs_i_1;
input  n_rst_c;
input  sck_33_c;
output vd_done;

    wire sig_prev_i, sig_prev_net_1, sig_old_i_0, GND, VCC;
    
    NOR2B sig_old_RNIERFT (.A(sig_prev_net_1), .B(sig_old_i_0), .Y(
        vd_done));
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(sck_33_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev (.D(cs_i_1), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        sig_prev_net_1));
    INV sig_old_RNO (.A(sig_prev_net_1), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module spi_ctl_12s_3_0(
       n_rst_c,
       sck_33_c,
       N_29,
       cs_i_1,
       cs_i_1_i
    );
input  n_rst_c;
input  sck_33_c;
output N_29;
output cs_i_1;
output cs_i_1_i;

    wire cnt_m1_0_a2_0, \cnt[14]_net_1 , \cnt[13]_net_1 , 
        cnt_m6_0_a2_6, cnt_m6_0_a2_0, \cnt[3]_net_1 , cnt_m5_0_a2_2, 
        cnt_m6_0_a2_2, \cnt[7]_net_1 , \cnt[8]_net_1 , \cnt[11]_net_1 , 
        \cnt[10]_net_1 , cnt_m7_0_a2_4, \cnt[5]_net_1 , cnt_m7_0_a2_3, 
        \cnt[6]_net_1 , cnt_m7_0_a2_1, \cnt[9]_net_1 , 
        state_tr0_0_a3_12, state_tr0_0_a3_6, state_tr0_0_a3_9, N_103, 
        \cnt[4]_net_1 , state_tr0_0_a3_8, state_tr0_0_a3_4, 
        state_tr0_0_a3_7, state_tr0_0_a3_2, \cnt[0]_net_1 , 
        \cnt[1]_net_1 , state_tr0_0_a3_1, \cnt[15]_net_1 , 
        \cnt[12]_net_1 , vd_stp_en_i_a3_9, vd_stp_en_i_a3_4, 
        vd_stp_en_i_a3_3, N_73, vd_stp_en_i_a3_8, vd_stp_en_i_a3_2, 
        vd_stp_en_i_a3_5, cnt_m6_0_a2_5_6, cnt_m6_0_a2_5_0, 
        cnt_m6_0_a2_5, \cnt[2]_net_1 , cnt_m5_0_a2_3, cnt_m2_0_a2_0, 
        cnt_m5_0_a2_1, cnt_m2_0_a2_2, cnt_m2_0_a2_1, N_74, 
        cnt_N_13_mux, N_33, N_31, cnt_N_7_mux_0_0, cnt_N_3_mux_0, 
        cnt_N_11_mux_2, cnt_N_15_mux, cnt_N_13_mux_0, N_30, 
        \state_RNO_4[0]_net_1 , N_26, N_24, N_22, N_20, N_97, N_18, 
        N_14, N_12, N_36, \cnt_RNO_0[6]_net_1 , cnt_n10, d_N_3_mux_1, 
        \cnt_RNO_1_1[10] , cnt_n0, cnt_n15, cnt_n14, cnt_n13, N_72, 
        cnt_n12, cnt_n11, cnt_n9, N_38, GND, VCC;
    
    NOR2B \cnt_RNO_2[6]  (.A(\cnt[4]_net_1 ), .B(\cnt[3]_net_1 ), .Y(
        cnt_m2_0_a2_2));
    XA1A \cnt_RNO[8]  (.A(\cnt[8]_net_1 ), .B(N_36), .C(cs_i_1), .Y(
        N_12));
    NOR2B \cnt_RNID4KA_0[1]  (.A(\cnt[1]_net_1 ), .B(\cnt[0]_net_1 ), 
        .Y(cnt_m2_0_a2_0));
    NOR3C \cnt_RNO_3[10]  (.A(\cnt[3]_net_1 ), .B(\cnt[5]_net_1 ), .C(
        cs_i_1), .Y(cnt_m7_0_a2_4));
    NOR3A \state_RNO_0[0]  (.A(state_tr0_0_a3_4), .B(\cnt[6]_net_1 ), 
        .C(\cnt[7]_net_1 ), .Y(state_tr0_0_a3_8));
    NOR3C \cnt_RNIM59L[9]  (.A(\cnt[9]_net_1 ), .B(\cnt[6]_net_1 ), .C(
        cnt_m6_0_a2_2), .Y(cnt_m6_0_a2_5));
    XA1A \cnt_RNO[2]  (.A(N_30), .B(\cnt[2]_net_1 ), .C(cs_i_1), .Y(
        N_24));
    DFN1C0 \cnt[2]  (.D(N_24), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[2]_net_1 ));
    DFN1C0 \cnt[8]  (.D(N_12), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[8]_net_1 ));
    DFN1C0 \cnt[1]  (.D(N_26), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[1]_net_1 ));
    OA1C \cnt_RNO_0[4]  (.A(\cnt[3]_net_1 ), .B(N_31), .C(
        \cnt[4]_net_1 ), .Y(N_97));
    DFN1C0 \cnt[11]  (.D(cnt_n11), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[11]_net_1 ));
    NOR3C \cnt_RNO_0[6]  (.A(cnt_m2_0_a2_1), .B(cnt_m2_0_a2_0), .C(
        cnt_m2_0_a2_2), .Y(cnt_N_7_mux_0_0));
    NOR2 \cnt_RNII0NU[11]  (.A(\cnt[11]_net_1 ), .B(\cnt[13]_net_1 ), 
        .Y(state_tr0_0_a3_1));
    NOR2B \cnt_RNO_1[15]  (.A(\cnt[14]_net_1 ), .B(\cnt[13]_net_1 ), 
        .Y(cnt_m1_0_a2_0));
    XA1A \cnt_RNO[3]  (.A(N_31), .B(\cnt[3]_net_1 ), .C(cs_i_1), .Y(
        N_22));
    OR2B \cnt_RNO_0[13]  (.A(cnt_N_13_mux), .B(\cnt[12]_net_1 ), .Y(
        N_72));
    NOR2B \cnt_RNILCKA[5]  (.A(\cnt[4]_net_1 ), .B(\cnt[5]_net_1 ), .Y(
        cnt_m5_0_a2_2));
    NOR3B \cnt_RNIOSSJ2[3]  (.A(cnt_m6_0_a2_6), .B(cnt_m6_0_a2_5), .C(
        N_31), .Y(cnt_N_13_mux));
    NOR3 \cnt_RNIIC141[15]  (.A(\cnt[14]_net_1 ), .B(\cnt[15]_net_1 ), 
        .C(\cnt[5]_net_1 ), .Y(vd_stp_en_i_a3_5));
    NOR3B \state_RNO_6[0]  (.A(\cnt[5]_net_1 ), .B(N_103), .C(
        \cnt[4]_net_1 ), .Y(state_tr0_0_a3_9));
    VCC VCC_i (.Y(VCC));
    NOR2 \cnt_RNIGUMU[10]  (.A(\cnt[10]_net_1 ), .B(\cnt[12]_net_1 ), 
        .Y(vd_stp_en_i_a3_2));
    INV \state_RNIIODF[0]  (.A(cs_i_1), .Y(cs_i_1_i));
    XA1 \cnt_RNO[1]  (.A(\cnt[0]_net_1 ), .B(\cnt[1]_net_1 ), .C(
        cs_i_1), .Y(N_26));
    NOR2B \cnt_RNIKBKA[2]  (.A(\cnt[2]_net_1 ), .B(\cnt[6]_net_1 ), .Y(
        cnt_m5_0_a2_1));
    DFN1C0 \cnt[6]  (.D(\cnt_RNO_0[6]_net_1 ), .CLK(sck_33_c), .CLR(
        n_rst_c), .Q(\cnt[6]_net_1 ));
    NOR3C \cnt_RNO_0[15]  (.A(cnt_m1_0_a2_0), .B(\cnt[12]_net_1 ), .C(
        cnt_N_13_mux), .Y(cnt_N_3_mux_0));
    OR2A \cnt_RNIBEUF[4]  (.A(\cnt[4]_net_1 ), .B(N_103), .Y(N_73));
    NOR3A \state_RNO_1[0]  (.A(state_tr0_0_a3_2), .B(\cnt[0]_net_1 ), 
        .C(\cnt[1]_net_1 ), .Y(state_tr0_0_a3_7));
    DFN1C0 \cnt[4]  (.D(N_20), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[4]_net_1 ));
    DFN1C0 \cnt[9]  (.D(cnt_n9), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[9]_net_1 ));
    NOR2A \cnt_RNO[0]  (.A(cs_i_1), .B(\cnt[0]_net_1 ), .Y(cnt_n0));
    OR3C \cnt_RNO_0[14]  (.A(\cnt[12]_net_1 ), .B(\cnt[13]_net_1 ), .C(
        cnt_N_13_mux), .Y(N_74));
    DFN1C0 \cnt[0]  (.D(cnt_n0), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[0]_net_1 ));
    NOR3B \cnt_RNO[4]  (.A(N_33), .B(cs_i_1), .C(N_97), .Y(N_20));
    OR3B \cnt_RNIOIIQ[4]  (.A(\cnt[3]_net_1 ), .B(\cnt[4]_net_1 ), .C(
        N_31), .Y(N_33));
    NOR2 \state_RNO_4[0]  (.A(\cnt[10]_net_1 ), .B(\cnt[8]_net_1 ), .Y(
        state_tr0_0_a3_2));
    DFN1C0 \state[0]  (.D(\state_RNO_4[0]_net_1 ), .CLK(sck_33_c), 
        .CLR(n_rst_c), .Q(cs_i_1));
    XA1 \cnt_RNO[6]  (.A(cnt_N_7_mux_0_0), .B(\cnt[6]_net_1 ), .C(
        cs_i_1), .Y(\cnt_RNO_0[6]_net_1 ));
    OR2B \cnt_RNICAHA1[7]  (.A(cnt_N_11_mux_2), .B(\cnt[7]_net_1 ), .Y(
        N_36));
    XA1 \cnt_RNO[15]  (.A(\cnt[15]_net_1 ), .B(cnt_N_3_mux_0), .C(
        cs_i_1), .Y(cnt_n15));
    XA1A \cnt_RNO[9]  (.A(\cnt[9]_net_1 ), .B(N_38), .C(cs_i_1), .Y(
        cnt_n9));
    GND GND_i (.Y(GND));
    NOR2B \cnt_RNO_5[10]  (.A(\cnt[8]_net_1 ), .B(\cnt[9]_net_1 ), .Y(
        cnt_m7_0_a2_1));
    NOR2 \cnt_RNIH8KA[2]  (.A(\cnt[3]_net_1 ), .B(\cnt[2]_net_1 ), .Y(
        N_103));
    OR2B \cnt_RNID4KA[1]  (.A(\cnt[1]_net_1 ), .B(\cnt[0]_net_1 ), .Y(
        N_30));
    DFN1C0 \cnt[13]  (.D(cnt_n13), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[13]_net_1 ));
    NOR3A \state_RNO_5[0]  (.A(state_tr0_0_a3_1), .B(\cnt[14]_net_1 ), 
        .C(\cnt[15]_net_1 ), .Y(state_tr0_0_a3_6));
    OR2A \cnt_RNO_0[9]  (.A(\cnt[8]_net_1 ), .B(N_36), .Y(N_38));
    DFN1C0 \cnt[7]  (.D(N_14), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[7]_net_1 ));
    NOR3C \state_RNO_2[0]  (.A(state_tr0_0_a3_6), .B(cs_i_1), .C(
        state_tr0_0_a3_9), .Y(state_tr0_0_a3_12));
    NOR3C \cnt_RNIF1751[2]  (.A(cnt_m5_0_a2_2), .B(cnt_m5_0_a2_1), .C(
        cnt_m5_0_a2_3), .Y(cnt_N_11_mux_2));
    DFN1C0 \cnt[10]  (.D(cnt_n10), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[10]_net_1 ));
    NOR3C \cnt_RNO_1[11]  (.A(cnt_m6_0_a2_5_0), .B(\cnt[3]_net_1 ), .C(
        cnt_m5_0_a2_2), .Y(cnt_m6_0_a2_5_6));
    XA1A \cnt_RNO[5]  (.A(\cnt[5]_net_1 ), .B(N_33), .C(cs_i_1), .Y(
        N_18));
    NOR2B \cnt_RNI69UF[3]  (.A(\cnt[3]_net_1 ), .B(cnt_m2_0_a2_0), .Y(
        cnt_m5_0_a2_3));
    NOR3C \cnt_RNI1K751[4]  (.A(vd_stp_en_i_a3_4), .B(vd_stp_en_i_a3_3)
        , .C(N_73), .Y(vd_stp_en_i_a3_9));
    DFN1C0 \cnt[3]  (.D(N_22), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[3]_net_1 ));
    NOR2B \cnt_RNO_2[11]  (.A(\cnt[10]_net_1 ), .B(\cnt[2]_net_1 ), .Y(
        cnt_m6_0_a2_5_0));
    XA1A \cnt_RNO[14]  (.A(\cnt[14]_net_1 ), .B(N_74), .C(cs_i_1), .Y(
        cnt_n14));
    NOR3C \cnt_RNIKBF13[10]  (.A(vd_stp_en_i_a3_2), .B(
        state_tr0_0_a3_1), .C(vd_stp_en_i_a3_5), .Y(vd_stp_en_i_a3_8));
    XNOR2 \cnt_RNO_1[10]  (.A(\cnt[10]_net_1 ), .B(\cnt[4]_net_1 ), .Y(
        \cnt_RNO_1_1[10] ));
    NOR3C \cnt_RNO_4[10]  (.A(\cnt[7]_net_1 ), .B(\cnt[6]_net_1 ), .C(
        cnt_m7_0_a2_1), .Y(cnt_m7_0_a2_3));
    OR2A \cnt_RNI58UF[2]  (.A(\cnt[2]_net_1 ), .B(N_30), .Y(N_31));
    NOR3B \cnt_RNO_0[11]  (.A(cnt_m6_0_a2_5), .B(cnt_m6_0_a2_5_6), .C(
        N_30), .Y(cnt_N_13_mux_0));
    NOR2 \cnt_RNISJKA[9]  (.A(\cnt[9]_net_1 ), .B(\cnt[7]_net_1 ), .Y(
        vd_stp_en_i_a3_4));
    XA1 \cnt_RNO[11]  (.A(\cnt[11]_net_1 ), .B(cnt_N_13_mux_0), .C(
        cs_i_1), .Y(cnt_n11));
    NOR2B \cnt_RNIFTMU[11]  (.A(\cnt[11]_net_1 ), .B(\cnt[10]_net_1 ), 
        .Y(cnt_m6_0_a2_0));
    NOR2 \cnt_RNIQHKA[6]  (.A(\cnt[8]_net_1 ), .B(\cnt[6]_net_1 ), .Y(
        vd_stp_en_i_a3_3));
    NOR3B \cnt_RNO_2[10]  (.A(cnt_m7_0_a2_4), .B(cnt_m7_0_a2_3), .C(
        N_31), .Y(cnt_N_15_mux));
    OR3C \state_RNO[0]  (.A(state_tr0_0_a3_8), .B(state_tr0_0_a3_7), 
        .C(state_tr0_0_a3_12), .Y(\state_RNO_4[0]_net_1 ));
    MX2B \cnt_RNO[10]  (.A(d_N_3_mux_1), .B(\cnt_RNO_1_1[10] ), .S(
        cnt_N_15_mux), .Y(cnt_n10));
    DFN1C0 \cnt[15]  (.D(cnt_n15), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[15]_net_1 ));
    AO1B \state_RNI7O4M4[0]  (.A(vd_stp_en_i_a3_9), .B(
        vd_stp_en_i_a3_8), .C(cs_i_1), .Y(N_29));
    NOR2B \cnt_RNO_1[6]  (.A(\cnt[2]_net_1 ), .B(\cnt[5]_net_1 ), .Y(
        cnt_m2_0_a2_1));
    NOR3C \cnt_RNITELE1[3]  (.A(cnt_m6_0_a2_0), .B(\cnt[3]_net_1 ), .C(
        cnt_m5_0_a2_2), .Y(cnt_m6_0_a2_6));
    NOR2B \cnt_RNIRIKA[7]  (.A(\cnt[7]_net_1 ), .B(\cnt[8]_net_1 ), .Y(
        cnt_m6_0_a2_2));
    NOR2B \cnt_RNO_0[10]  (.A(\cnt[10]_net_1 ), .B(cs_i_1), .Y(
        d_N_3_mux_1));
    NOR2 \state_RNO_3[0]  (.A(\cnt[9]_net_1 ), .B(\cnt[12]_net_1 ), .Y(
        state_tr0_0_a3_4));
    DFN1C0 \cnt[5]  (.D(N_18), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[5]_net_1 ));
    XA1A \cnt_RNO[13]  (.A(\cnt[13]_net_1 ), .B(N_72), .C(cs_i_1), .Y(
        cnt_n13));
    XA1 \cnt_RNO[12]  (.A(\cnt[12]_net_1 ), .B(cnt_N_13_mux), .C(
        cs_i_1), .Y(cnt_n12));
    DFN1C0 \cnt[12]  (.D(cnt_n12), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[12]_net_1 ));
    XA1 \cnt_RNO[7]  (.A(\cnt[7]_net_1 ), .B(cnt_N_11_mux_2), .C(
        cs_i_1), .Y(N_14));
    DFN1C0 \cnt[14]  (.D(cnt_n14), .CLK(sck_33_c), .CLR(n_rst_c), .Q(
        \cnt[14]_net_1 ));
    
endmodule


module spi_rx_12s_3_0(
       cur_vd,
       vd_done,
       cs_i_1_i,
       sck_33_c,
       n_rst_c,
       din_fb_c
    );
output [11:0] cur_vd;
output vd_done;
output cs_i_1_i;
input  sck_33_c;
input  n_rst_c;
input  din_fb_c;

    wire N_29, cs_i_1, GND, VCC;
    
    spi_stp_12s_1_6_0 VD_STP (.cur_vd({cur_vd[11], cur_vd[10], 
        cur_vd[9], cur_vd[8], cur_vd[7], cur_vd[6], cur_vd[5], 
        cur_vd[4], cur_vd[3], cur_vd[2], cur_vd[1], cur_vd[0]}), .N_29(
        N_29), .din_fb_c(din_fb_c), .n_rst_c(n_rst_c), .sck_33_c(
        sck_33_c));
    sig_gen_0_0 SPI_RDYSIG (.cs_i_1(cs_i_1), .n_rst_c(n_rst_c), 
        .sck_33_c(sck_33_c), .vd_done(vd_done));
    VCC VCC_i (.Y(VCC));
    spi_ctl_12s_3_0 SPICTL (.n_rst_c(n_rst_c), .sck_33_c(sck_33_c), 
        .N_29(N_29), .cs_i_1(cs_i_1), .cs_i_1_i(cs_i_1_i));
    GND GND_i (.Y(GND));
    
endmodule


module integral_calc_13s_0_4_1(
       sr_old,
       sr_new,
       sr_new_0_0,
       sr_new_1_0,
       integral,
       sr_old_0_0,
       integral_i,
       integral_0_0,
       integral_1_0,
       calc_int,
       int_done,
       n_rst_c,
       clk_c
    );
input  [12:0] sr_old;
input  [12:0] sr_new;
input  sr_new_0_0;
input  sr_new_1_0;
output [25:6] integral;
input  sr_old_0_0;
output [25:24] integral_i;
output integral_0_0;
output integral_1_0;
input  calc_int;
output int_done;
input  n_rst_c;
input  clk_c;

    wire \un1_integ[25] , \un1_next_int_0_iv_0[13] , 
        next_int_0_sqmuxa_1, next_int_1_sqmuxa, int_done_0, 
        \state[1]_net_1 , \state[0]_net_1 , N_12, N_10, 
        \DWACT_FINC_E[0] , N_5, \DWACT_FINC_E[4] , N_2, 
        \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , N_12_0, N_10_0, 
        \DWACT_FINC_E_0[0] , N_5_0, \DWACT_FINC_E_0[4] , N_2_0, 
        \DWACT_FINC_E_0[7] , \DWACT_FINC_E_0[6] , 
        ADD_26x26_fast_I254_Y_0, \un1_next_int_0_iv[13] , 
        ADD_26x26_fast_I255_Y_0, ADD_26x26_fast_I253_Y_0, 
        ADD_26x26_fast_I252_Y_0, ADD_26x26_fast_I249_Y_0, 
        ADD_26x26_fast_I248_Y_0, ADD_26x26_fast_I246_Y_0, 
        ADD_26x26_fast_I247_Y_0, ADD_26x26_fast_I204_Y_3, N517, N502, 
        ADD_26x26_fast_I204_Y_2, N398, ADD_26x26_fast_I204_Y_0, N455, 
        ADD_26x26_fast_I205_Y_3, N504, N519, ADD_26x26_fast_I205_Y_2, 
        N400, ADD_26x26_fast_I205_Y_0, N457, ADD_26x26_fast_I251_Y_0, 
        ADD_26x26_fast_I250_Y_0, ADD_26x26_fast_I207_Y_2, 
        ADD_26x26_fast_I207_un1_Y_0, N524, ADD_26x26_fast_I207_Y_1, 
        N404, N461, ADD_26x26_fast_I206_Y_2, 
        ADD_26x26_fast_I206_un1_Y_0, N522, ADD_26x26_fast_I206_Y_1, 
        N459, N452, ADD_26x26_fast_I206_Y_0, N399, N402, 
        ADD_26x26_fast_I244_Y_0, ADD_26x26_fast_I245_Y_0, 
        ADD_26x26_fast_I210_Y_1, N529, N514, ADD_26x26_fast_I210_Y_0, 
        I136_un1_Y, ADD_26x26_fast_I211_Y_1, N516, N531, 
        ADD_26x26_fast_I211_Y_0, N469, N462, ADD_26x26_fast_I212_Y_0, 
        N533, N518, ADD_26x26_fast_I213_Y_0, N535, N520, 
        ADD_26x26_fast_I243_Y_0, ADD_26x26_fast_I241_Y_0, 
        \state_RNIJ1O9E[0]_net_1 , ADD_26x26_fast_I242_Y_0, 
        \un1_next_int[12] , ADD_26x26_fast_I240_Y_0, 
        \state_RNI00AMD[0]_net_1 , ADD_26x26_fast_I209_Y_1, 
        ADD_26x26_fast_I209_un1_Y_0, N528, ADD_26x26_fast_I209_Y_0, 
        N465, N458, ADD_26x26_fast_I208_Y_1, 
        ADD_26x26_fast_I208_un1_Y_0, N526, ADD_26x26_fast_I208_Y_0, 
        N456, N463, ADD_26x26_fast_I204_un1_Y_0, 
        ADD_26x26_fast_I239_Y_0, \state_RNISE23D[0]_net_1 , 
        ADD_26x26_fast_I212_un1_Y_0, N480, N488, N442, N483, 
        I160_un1_Y, N506, N485, I161_un1_Y, N508, N487, I162_un1_Y, 
        N510, N489, I163_un1_Y, N512, ADD_26x26_fast_I237_Y_0, 
        \state_RNIU2U5B[0]_net_1 , ADD_26x26_fast_I235_Y_0, 
        \un2_next_int_m[5] , \un1_next_int_iv_1[5] , \integ[5]_net_1 , 
        ADD_26x26_fast_I236_Y_0, \un1_next_int[6] , 
        ADD_26x26_fast_I234_Y_0, \integ[4]_net_1 , \un1_next_int[4] , 
        ADD_26x26_fast_I232_Y_0, \integ[2]_net_1 , \un1_next_int[2] , 
        ADD_26x26_fast_I127_Y_0, ADD_26x26_fast_I125_Y_0, 
        ADD_26x26_fast_I231_Y_0, \integ[1]_net_1 , \un1_next_int[1] , 
        \un1_next_int_iv_0[10] , \inf_abs1[10]_net_1 , 
        \un1_next_int_iv_0[11] , \inf_abs1[11]_net_1 , 
        \un1_next_int_iv_1[9] , \un1_next_int_iv_0[9] , 
        \inf_abs0_m[9] , \inf_abs1[9]_net_1 , \un1_next_int_iv_1[7] , 
        \un1_next_int_iv_0[7] , \inf_abs0_m[7] , \inf_abs1[7]_net_1 , 
        \un1_next_int_iv_0[4] , \inf_abs1[4]_net_1 , 
        \un1_next_int_iv_0[6] , \inf_abs1[6]_net_1 , 
        ADD_26x26_fast_I230_Y_0, \integ[0]_net_1 , N_3, 
        \un1_next_int_iv_0[12] , \inf_abs1_a_1[12] , 
        \un1_next_int_iv_1[0] , \un18_next_int_m[0] , \inf_abs1_m[0] , 
        \un2_next_int_m[0] , \inf_abs0_m[5] , \un18_next_int_m[5] , 
        \inf_abs1_m[5] , \un1_next_int_iv_1[8] , \inf_abs0_m[8] , 
        \un18_next_int_m[8] , \inf_abs1_m[8] , \un1_next_int_iv_0[3] , 
        \inf_abs1[3]_net_1 , \un1_next_int_iv_0[2] , 
        \inf_abs1[2]_net_1 , \un1_next_int_iv_1[1] , 
        \un18_next_int_m[1] , \inf_abs1_m[1] , \un2_next_int_m[1] , 
        \inf_abs0_m[1] , \un2_next_int_m[12] , 
        \state_RNIJL492[0]_net_1 , \inf_abs0_m[0] , \un1_next_int[8] , 
        \un2_next_int_m[8] , \un1_integ[0] , \inf_abs0_m[4] , 
        \un2_next_int_m[4] , \inf_abs0_m[6] , \un2_next_int_m[6] , 
        \un2_next_int_m[7] , \inf_abs0_m[10] , \un2_next_int_m[10] , 
        \inf_abs0_m[11] , \un2_next_int_m[11] , \un1_integ[3] , 
        \un1_next_int[3] , \integ[3]_net_1 , N491, I204_un1_Y, 
        I194_un1_Y, \un1_integ[9] , \un1_integ[13] , N525, I190_un1_Y, 
        \un1_integ[12] , N527, I191_un1_Y, \un1_integ[21] , I176_un1_Y, 
        \un1_integ[5] , \un1_integ[1] , \un1_integ[17] , I212_un1_Y, 
        \un1_integ[15] , N521, I188_un1_Y, \un1_integ[23] , I172_un1_Y, 
        \un1_integ[20] , I178_un1_Y, N405, N401, I205_un1_Y, N658, 
        I211_un1_Y, N493, N532, \un1_integ[22] , I174_un1_Y, 
        \un1_integ[18] , \un1_integ[24] , \un1_integ[14] , N523, 
        I189_un1_Y, \un1_integ[6] , \un1_integ[8] , I213_un1_Y, N536, 
        \un1_integ[2] , \un1_integ[16] , \un1_integ[7] , 
        \un1_integ[19] , I210_un1_Y, \un1_integ[10] , I193_un1_Y, 
        \un1_integ[11] , I192_un1_Y, \un1_integ[4] , 
        \un2_next_int_m[9] , N530, \inf_abs0_m[3] , 
        \un2_next_int_m[3] , \inf_abs0_m[2] , \un2_next_int_m[2] , 
        \inf_abs1_a_1[2] , \inf_abs0[2]_net_1 , \inf_abs0_a_0[2] , 
        \inf_abs1_a_1[3] , \inf_abs0[3]_net_1 , \inf_abs0_a_0[3] , 
        N467, N460, N468, \inf_abs0[9]_net_1 , \inf_abs0_a_0[9] , 
        \inf_abs1_a_1[9] , I96_un1_Y, N414, N324, N323, I195_un1_Y, 
        N408, I90_un1_Y, N411, N410, N409, N413, N403, N407, N478, 
        N477, N406, N470, I146_un1_Y, N466, \state_RNO_3[0] , N473, 
        I158_un1_Y, N482, N481, N490, N479, I108_un1_Y, N426, N338, 
        N342, N341, N430, N427, N339, N431, N333, N336, N424, N421, 
        N420, N347, N351, N350, N348, N474, N425, N345, N429, N472, 
        N423, N419, N354, N433, N330, N432, N428, N335, N332, N415, 
        N471, N422, N418, N475, N476, N434, N484, N326, N329, 
        I50_un1_Y, N353, N344, N436, \inf_abs0[4]_net_1 , 
        \inf_abs0[6]_net_1 , \inf_abs0[7]_net_1 , \inf_abs0[10]_net_1 , 
        \inf_abs0[11]_net_1 , \inf_abs0_a_0[4] , \inf_abs0_a_0[6] , 
        \inf_abs0_a_0[7] , \inf_abs0_a_0[10] , \inf_abs0_a_0[11] , 
        \inf_abs1_a_1[4] , \inf_abs1_a_1[6] , \inf_abs1_a_1[7] , 
        \inf_abs1_a_1[10] , \inf_abs1_a_1[11] , N417, N416, N486, N439, 
        N321, N327, N437, N318, N438, N320, N317, N464, I148_un1_Y, 
        \state_RNO_4[1] , I121_un1_Y, N440, N441, N435, I74_un1_Y, 
        I118_un1_Y, I150_un1_Y, \inf_abs0_a_0[8] , \inf_abs1_a_1[8] , 
        \inf_abs0_a_0[5] , \inf_abs1_a_1[5] , \inf_abs0_a_0[12] , 
        \inf_abs0_a_0[1] , \inf_abs1_a_1[1] , N_3_0, \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[5] , N_4, \DWACT_FINC_E[3] , N_6, N_7, N_8, 
        \DWACT_FINC_E[1] , N_9, N_11, N_3_1, \DWACT_FINC_E_0[2] , 
        \DWACT_FINC_E_0[5] , N_4_0, \DWACT_FINC_E_0[3] , N_6_0, N_7_0, 
        N_8_0, \DWACT_FINC_E_0[1] , N_9_0, N_11_0, GND, VCC;
    
    AO1 un1_integ_0_0_ADD_26x26_fast_I56_Y (.A(N341), .B(N345), .C(
        N344), .Y(N424));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I148_un1_Y (.A(N479), .B(N472), 
        .Y(I148_un1_Y));
    NOR2 inf_abs1_a_1_I_15 (.A(sr_old[3]), .B(sr_old[4]), .Y(
        \DWACT_FINC_E[1] ));
    XNOR2 inf_abs1_a_1_I_23 (.A(sr_old[8]), .B(N_6), .Y(
        \inf_abs1_a_1[8] ));
    DFN1C0 \state[0]  (.D(\state_RNO_3[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[0]_net_1 ));
    XNOR2 inf_abs1_a_1_I_17 (.A(sr_old[6]), .B(N_8), .Y(
        \inf_abs1_a_1[6] ));
    DFN1E0C0 \integ[13]  (.D(\un1_integ[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[13]));
    DFN1E0C0 \integ[24]  (.D(\un1_integ[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[24]));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I245_Y_0 (.A(integral[15]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I245_Y_0));
    OR2 \state_RNI42RG[1]  (.A(next_int_0_sqmuxa_1), .B(
        next_int_1_sqmuxa), .Y(\un1_next_int_0_iv_0[13] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I61_Y (.A(N336), .B(N339), .Y(
        N429));
    NOR2B \state_RNIOJ2D[0]  (.A(sr_new[8]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[8] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I7_P0N (.A(integral[7]), .B(
        \state_RNIU2U5B[0]_net_1 ), .Y(N339));
    NOR3B inf_abs0_a_0_I_19 (.A(\DWACT_FINC_E_0[2] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[6]), .Y(N_7_0));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I248_Y_0 (.A(integral[18]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I248_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I172_un1_Y (.A(N521), .B(N506), 
        .Y(I172_un1_Y));
    NOR3B inf_abs0_a_0_I_16 (.A(\DWACT_FINC_E_0[1] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[5]), .Y(N_8_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I41_Y (.A(integral[16]), .B(
        integral[17]), .C(\un1_next_int_0_iv_0[13] ), .Y(N409));
    OA1 un1_integ_0_0_ADD_26x26_fast_I204_un1_Y (.A(N533), .B(
        I194_un1_Y), .C(ADD_26x26_fast_I204_un1_Y_0), .Y(I204_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I86_Y (.A(N404), .B(N408), .Y(
        N457));
    OR3 \state_RNIPR8F5[1]  (.A(\inf_abs0_m[8] ), .B(
        \un18_next_int_m[8] ), .C(\inf_abs1_m[8] ), .Y(
        \un1_next_int_iv_1[8] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I98_Y (.A(N420), .B(N417), .C(
        N416), .Y(N469));
    NOR2B \state_RNIIFGM3_0[0]  (.A(next_int_1_sqmuxa), .B(
        \inf_abs0[9]_net_1 ), .Y(\inf_abs0_m[9] ));
    NOR3A \state_RNIQ44M[1]  (.A(\state[1]_net_1 ), .B(sr_old_0_0), .C(
        sr_old[8]), .Y(\un18_next_int_m[8] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I176_un1_Y (.A(N525), .B(N510), 
        .Y(I176_un1_Y));
    OR3 \state_RNIK4AP1[0]  (.A(\un18_next_int_m[0] ), .B(
        \inf_abs1_m[0] ), .C(\un2_next_int_m[0] ), .Y(
        \un1_next_int_iv_1[0] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I158_un1_Y (.A(N489), .B(N482), 
        .Y(I158_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I150_un1_Y (.A(N481), .B(N474), 
        .Y(I150_un1_Y));
    XA1A \state_RNIRD0C6[1]  (.A(sr_old[12]), .B(\inf_abs1[11]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[11] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I51_Y (.A(N354), .B(N351), .Y(
        N419));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y (.A(
        ADD_26x26_fast_I230_Y_0), .B(\state_RNIJL492[0]_net_1 ), .Y(
        \un1_integ[0] ));
    NOR2B inf_abs1_a_1_I_34 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .Y(N_2_0));
    NOR2B \state_RNI851A1[1]  (.A(\inf_abs1_a_1[1] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[1] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I253_Y (.A(I172_un1_Y), .B(
        ADD_26x26_fast_I206_Y_2), .C(ADD_26x26_fast_I253_Y_0), .Y(
        \un1_integ[23] ));
    DFN1E0C0 \integ[21]  (.D(\un1_integ[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[21]));
    XNOR2 inf_abs1_a_1_I_7 (.A(sr_old[2]), .B(N_12_0), .Y(
        \inf_abs1_a_1[2] ));
    DFN1E0C0 \integ_1[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done), .Q(integral_1_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I190_un1_Y (.A(N487), .B(
        I162_un1_Y), .C(N526), .Y(I190_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I146_Y (.A(I146_un1_Y), .B(N469), 
        .Y(N523));
    AO1 un1_integ_0_0_ADD_26x26_fast_I142_Y (.A(N473), .B(N466), .C(
        N465), .Y(N519));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I244_Y_0 (.A(integral[14]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I244_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I231_Y (.A(
        ADD_26x26_fast_I231_Y_0), .B(N442), .Y(\un1_integ[1] ));
    AND3 inf_abs1_a_1_I_24 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E_0[4] ));
    XNOR2 inf_abs1_a_1_I_32 (.A(sr_old[11]), .B(N_3_0), .Y(
        \inf_abs1_a_1[11] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I155_Y (.A(N486), .B(N478), .Y(
        N532));
    DFN1E0C0 \integ[15]  (.D(\un1_integ[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[15]));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I213_un1_Y (.A(N536), .B(
        \state_RNIJL492[0]_net_1 ), .C(N520), .Y(I213_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I103_Y (.A(N421), .B(N425), .Y(
        N474));
    XA1A \state_RNICL3K4[1]  (.A(sr_old_0_0), .B(\inf_abs1[7]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[7] ));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I125_Y (.A(N399), .B(
        ADD_26x26_fast_I125_Y_0), .C(N456), .Y(N502));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_1 (.A(
        ADD_26x26_fast_I209_un1_Y_0), .B(N528), .C(
        ADD_26x26_fast_I209_Y_0), .Y(ADD_26x26_fast_I209_Y_1));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I97_Y (.A(N415), .B(N419), .Y(
        N468));
    NOR3A \state_RNIIS3M_0[1]  (.A(\state[1]_net_1 ), .B(sr_old_0_0), 
        .C(sr_old[0]), .Y(\un18_next_int_m[0] ));
    NOR2A \state_RNI5SP2[0]  (.A(\state[0]_net_1 ), .B(sr_new[12]), .Y(
        next_int_1_sqmuxa));
    AO1 un1_integ_0_0_ADD_26x26_fast_I94_Y (.A(N416), .B(N413), .C(
        I90_un1_Y), .Y(N465));
    NOR2 inf_abs0_a_0_I_6 (.A(sr_new[0]), .B(sr_new[1]), .Y(N_12));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I81_Y (.A(N399), .B(N403), .Y(
        N452));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I151_Y (.A(N474), .B(N482), .Y(
        N528));
    AND3 inf_abs1_a_1_I_22 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_6));
    OR2 un1_integ_0_0_ADD_26x26_fast_I74_Y (.A(I74_un1_Y), .B(N317), 
        .Y(N442));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I238_Y (.A(\un1_next_int[8] ), 
        .B(integral[8]), .C(N658), .Y(\un1_integ[8] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I121_Y (.A(I121_un1_Y), .B(N440), 
        .Y(N493));
    NOR3B \state_RNIM7D02[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[5] ), .Y(\un2_next_int_m[5] ));
    NOR3 inf_abs0_a_0_I_10 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2])
        , .Y(\DWACT_FINC_E[0] ));
    NOR3B \state_RNI333A2[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[4]_net_1 ), .Y(\un2_next_int_m[4] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I5_P0N (.A(\un2_next_int_m[5] ), 
        .B(\un1_next_int_iv_1[5] ), .C(\integ[5]_net_1 ), .Y(N333));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I236_Y_0 (.A(integral[6]), .B(
        \un1_next_int[6] ), .Y(ADD_26x26_fast_I236_Y_0));
    NOR3B \state_RNISRAN[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), .C(
        \inf_abs0_a_0[1] ), .Y(\un2_next_int_m[1] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I246_Y (.A(I213_un1_Y), .B(
        ADD_26x26_fast_I213_Y_0), .C(ADD_26x26_fast_I246_Y_0), .Y(
        \un1_integ[16] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I252_Y_0 (.A(integral[22]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I252_Y_0));
    NOR3B \state_RNIIFGM3[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[9]_net_1 ), .Y(\un2_next_int_m[9] ));
    MX2 \inf_abs0[6]  (.A(sr_new[6]), .B(\inf_abs0_a_0[6] ), .S(
        sr_new_1_0), .Y(\inf_abs0[6]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I39_Y (.A(integral[17]), .B(
        integral[18]), .C(\un1_next_int_0_iv_0[13] ), .Y(N407));
    OA1B un1_integ_0_0_ADD_26x26_fast_I32_Y (.A(integral[21]), .B(
        integral[20]), .C(\un1_next_int_0_iv_0[13] ), .Y(N400));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I194_un1_Y (.A(N480), .B(N488), 
        .C(N442), .Y(I194_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I108_un1_Y (.A(N430), .B(N427), 
        .Y(I108_un1_Y));
    NOR2A inf_abs0_a_0_I_11 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .Y(
        N_10));
    AO1B un1_integ_0_0_ADD_26x26_fast_I125_Y_0 (.A(integral[23]), .B(
        integral[24]), .C(\un1_next_int_0_iv_0[13] ), .Y(
        ADD_26x26_fast_I125_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I100_Y (.A(N422), .B(N419), .C(
        N418), .Y(N471));
    OR2 un1_integ_0_0_ADD_26x26_fast_I12_P0N (.A(integral[12]), .B(
        \un1_next_int[12] ), .Y(N354));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I10_G0N (.A(integral[10]), .B(
        \state_RNI00AMD[0]_net_1 ), .Y(N347));
    DFN1E0C0 \integ[12]  (.D(\un1_integ[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[12]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I109_Y (.A(N431), .B(N427), .Y(
        N480));
    XNOR2 inf_abs1_a_1_I_35 (.A(sr_old[12]), .B(N_2_0), .Y(
        \inf_abs1_a_1[12] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I205_Y_0 (.A(integral[22]), .B(
        integral[23]), .C(\un1_next_int_0_iv_0[13] ), .Y(
        ADD_26x26_fast_I205_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I115_Y (.A(N437), .B(N433), .Y(
        N486));
    NOR2B \state_RNI333A2_0[0]  (.A(\inf_abs0[4]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[4] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I12_G0N (.A(integral[12]), .B(
        \un1_next_int[12] ), .Y(N353));
    OR2 \state_RNIJL492[0]  (.A(\un1_next_int_iv_1[0] ), .B(
        \inf_abs0_m[0] ), .Y(\state_RNIJL492[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_0 (.A(N456), .B(N463), .C(
        N455), .Y(ADD_26x26_fast_I208_Y_0));
    INV \integ_RNIJ176[24]  (.A(integral[24]), .Y(integral_i[24]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I111_Y (.A(N433), .B(N429), .Y(
        N482));
    OR2 \state_RNI5S0T7[1]  (.A(\un1_next_int_iv_0[7] ), .B(
        \inf_abs0_m[7] ), .Y(\un1_next_int_iv_1[7] ));
    NOR2A inf_abs1_a_1_I_25 (.A(\DWACT_FINC_E_0[4] ), .B(sr_old[8]), 
        .Y(N_5_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I2_P0N (.A(\un1_next_int[2] ), .B(
        \integ[2]_net_1 ), .Y(N324));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I250_Y_0 (.A(integral[20]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I250_Y_0));
    OR2 \state_RNIAVHC9[1]  (.A(\un1_next_int_iv_0[9] ), .B(
        \inf_abs0_m[9] ), .Y(\un1_next_int_iv_1[9] ));
    NOR3A inf_abs1_a_1_I_27 (.A(\DWACT_FINC_E_0[4] ), .B(sr_old[8]), 
        .C(sr_old[9]), .Y(N_4));
    DFN1E0C0 \integ[10]  (.D(\un1_integ[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[10]));
    OA1 un1_integ_0_0_ADD_26x26_fast_I188_un1_Y (.A(N483), .B(
        I160_un1_Y), .C(N522), .Y(I188_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I6_G0N (.A(\un1_next_int[6] ), 
        .B(integral[6]), .Y(N335));
    MX2 \inf_abs1[10]  (.A(sr_old[10]), .B(\inf_abs1_a_1[10] ), .S(
        sr_old_0_0), .Y(\inf_abs1[10]_net_1 ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I249_Y (.A(I210_un1_Y), .B(
        ADD_26x26_fast_I210_Y_1), .C(ADD_26x26_fast_I249_Y_0), .Y(
        \un1_integ[19] ));
    GND GND_i (.Y(GND));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I146_un1_Y (.A(N477), .B(N470), 
        .Y(I146_un1_Y));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I246_Y_0 (.A(integral[16]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I246_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I6_P0N (.A(\un1_next_int[6] ), .B(
        integral[6]), .Y(N336));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I212_un1_Y_0 (.A(N480), .B(N488)
        , .C(N442), .Y(ADD_26x26_fast_I212_un1_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I1_G0N (.A(\integ[1]_net_1 ), 
        .B(\un1_next_int[1] ), .Y(N320));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I107_Y (.A(N425), .B(N429), .Y(
        N478));
    OR3 \state_RNIH89U7[0]  (.A(\inf_abs0_m[4] ), .B(
        \un1_next_int_iv_0[4] ), .C(\un2_next_int_m[4] ), .Y(
        \un1_next_int[4] ));
    XNOR2 inf_abs1_a_1_I_9 (.A(sr_old[3]), .B(N_11), .Y(
        \inf_abs1_a_1[3] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I38_Y (.A(integral[18]), .B(
        integral[17]), .C(\un1_next_int_0_iv_0[13] ), .Y(N406));
    OA1 un1_integ_0_0_ADD_26x26_fast_I209_un1_Y_0 (.A(N489), .B(
        I163_un1_Y), .C(N512), .Y(ADD_26x26_fast_I209_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_3 (.A(N504), .B(N519), .C(
        ADD_26x26_fast_I205_Y_2), .Y(ADD_26x26_fast_I205_Y_3));
    AX1D un1_integ_0_0_ADD_26x26_fast_I255_Y (.A(I204_un1_Y), .B(
        ADD_26x26_fast_I204_Y_3), .C(ADD_26x26_fast_I255_Y_0), .Y(
        \un1_integ[25] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I204_Y_0 (.A(integral[24]), .B(
        integral[23]), .C(\un1_next_int_0_iv_0[13] ), .Y(
        ADD_26x26_fast_I204_Y_0));
    MX2 \inf_abs0[4]  (.A(sr_new[4]), .B(\inf_abs0_a_0[4] ), .S(
        sr_new_1_0), .Y(\inf_abs0[4]_net_1 ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I243_Y (.A(N525), .B(I190_un1_Y), 
        .C(ADD_26x26_fast_I243_Y_0), .Y(\un1_integ[13] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I231_Y_0 (.A(\integ[1]_net_1 ), 
        .B(\un1_next_int[1] ), .Y(ADD_26x26_fast_I231_Y_0));
    OR2 \state_RNI8BI43[0]  (.A(\un1_next_int_iv_1[1] ), .B(
        \inf_abs0_m[1] ), .Y(\un1_next_int[1] ));
    OA1A \state_RNIMRU36[1]  (.A(sr_old[12]), .B(\inf_abs1_a_1[12] ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[12] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I69_Y (.A(N324), .B(N327), .Y(
        N437));
    AO1 un1_integ_0_0_ADD_26x26_fast_I62_Y (.A(N332), .B(N336), .C(
        N335), .Y(N430));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I193_un1_Y (.A(N532), .B(N493), 
        .Y(I193_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I153_Y (.A(N484), .B(N476), .Y(
        N530));
    OR2 \state_RNIU2U5B[0]  (.A(\un1_next_int_iv_1[7] ), .B(
        \un2_next_int_m[7] ), .Y(\state_RNIU2U5B[0]_net_1 ));
    NOR2B \state_RNI62LO3[0]  (.A(\inf_abs0[10]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[10] ));
    XNOR2 inf_abs0_a_0_I_7 (.A(sr_new[2]), .B(N_12), .Y(
        \inf_abs0_a_0[2] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I7_G0N (.A(integral[7]), .B(
        \state_RNIU2U5B[0]_net_1 ), .Y(N338));
    OA1A un1_integ_0_0_ADD_26x26_fast_I49_Y (.A(
        \un1_next_int_0_iv[13] ), .B(integral[13]), .C(N354), .Y(N417));
    OA1B un1_integ_0_0_ADD_26x26_fast_I42_Y (.A(integral[15]), .B(
        integral[16]), .C(\un1_next_int_0_iv_0[13] ), .Y(N410));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I145_Y (.A(N476), .B(N468), .Y(
        N522));
    OR3 \state_RNI73855[0]  (.A(\inf_abs0_m[2] ), .B(
        \un1_next_int_iv_0[2] ), .C(\un2_next_int_m[2] ), .Y(
        \un1_next_int[2] ));
    MX2 \inf_abs1[4]  (.A(sr_old[4]), .B(\inf_abs1_a_1[4] ), .S(
        sr_old[12]), .Y(\inf_abs1[4]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I10_P0N (.A(integral[10]), .B(
        \state_RNI00AMD[0]_net_1 ), .Y(N348));
    OR2 un1_integ_0_0_ADD_26x26_fast_I1_P0N (.A(\integ[1]_net_1 ), .B(
        \un1_next_int[1] ), .Y(N321));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I192_un1_Y (.A(N530), .B(N491), 
        .Y(I192_un1_Y));
    NOR3A inf_abs0_a_0_I_13 (.A(\DWACT_FINC_E[0] ), .B(sr_new[4]), .C(
        sr_new[3]), .Y(N_9_0));
    MX2 \inf_abs0[9]  (.A(sr_new[9]), .B(\inf_abs0_a_0[9] ), .S(
        sr_new[12]), .Y(\inf_abs0[9]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I141_Y (.A(N464), .B(N472), .Y(
        N518));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I93_Y (.A(N411), .B(N415), .Y(
        N464));
    AO1B un1_integ_0_0_ADD_26x26_fast_I37_Y (.A(integral[19]), .B(
        integral[18]), .C(\un1_next_int_0_iv_0[13] ), .Y(N405));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I0_G0N (.A(\integ[0]_net_1 ), 
        .B(N_3), .Y(N317));
    NOR3B \state_RNIVGQF[0]  (.A(\state[0]_net_1 ), .B(sr_new[0]), .C(
        sr_new_0_0), .Y(\inf_abs0_m[0] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I73_Y (.A(N318), .B(N321), .Y(
        N441));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I59_Y (.A(N342), .B(N339), .Y(
        N427));
    AO1 un1_integ_0_0_ADD_26x26_fast_I52_Y (.A(N347), .B(N351), .C(
        N350), .Y(N420));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I211_un1_Y (.A(N516), .B(N493), 
        .C(N532), .Y(I211_un1_Y));
    NOR2A \state_RNO[1]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 ), 
        .Y(\state_RNO_4[1] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I34_Y (.A(integral[19]), .B(
        integral[20]), .C(\un1_next_int_0_iv_0[13] ), .Y(N402));
    NOR3B \state_RNIKUA24[0]  (.A(sr_new_1_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[11]_net_1 ), .Y(\un2_next_int_m[11] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I236_Y (.A(N485), .B(I161_un1_Y), 
        .C(ADD_26x26_fast_I236_Y_0), .Y(\un1_integ[6] ));
    OR3 \state_RNICCC3A[0]  (.A(\inf_abs0_m[6] ), .B(
        \un1_next_int_iv_0[6] ), .C(\un2_next_int_m[6] ), .Y(
        \un1_next_int[6] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I150_Y (.A(I150_un1_Y), .B(N473), 
        .Y(N527));
    DFN1E0C0 \integ[0]  (.D(\un1_integ[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_done), .Q(\integ[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I120_Y (.A(N439), .B(N442), .C(
        N438), .Y(N491));
    AO1 un1_integ_0_0_ADD_26x26_fast_I104_Y (.A(N426), .B(N423), .C(
        N422), .Y(N475));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I159_Y (.A(N490), .B(N482), .Y(
        N536));
    NOR2B \state_RNI6G123[1]  (.A(\inf_abs1_a_1[5] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[5] ));
    VCC VCC_i (.Y(VCC));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I129_Y (.A(N460), .B(N452), .Y(
        N506));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I113_Y (.A(N435), .B(N431), .Y(
        N484));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I241_Y_0 (.A(integral[11]), .B(
        \state_RNIJ1O9E[0]_net_1 ), .Y(ADD_26x26_fast_I241_Y_0));
    XNOR2 inf_abs0_a_0_I_28 (.A(sr_new[10]), .B(N_4_0), .Y(
        \inf_abs0_a_0[10] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I89_Y (.A(N411), .B(N407), .Y(
        N460));
    AO1 un1_integ_0_0_ADD_26x26_fast_I68_Y (.A(N323), .B(N327), .C(
        N326), .Y(N436));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_0 (.A(N469), .B(N462), .C(
        N461), .Y(ADD_26x26_fast_I211_Y_0));
    NOR3A \state_RNIN14M[1]  (.A(\state[1]_net_1 ), .B(sr_old_0_0), .C(
        sr_old[5]), .Y(\un18_next_int_m[5] ));
    DFN1E0C0 \integ[4]  (.D(\un1_integ[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_done), .Q(\integ[4]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I108_Y (.A(I108_un1_Y), .B(N426), 
        .Y(N479));
    XA1A \state_RNIQQ2E2[1]  (.A(sr_old_0_0), .B(\inf_abs1[2]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[2] ));
    NOR3 inf_abs1_a_1_I_18 (.A(sr_old[4]), .B(sr_old[3]), .C(sr_old[5])
        , .Y(\DWACT_FINC_E[2] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I3_G0N (.A(\integ[3]_net_1 ), 
        .B(\un1_next_int[3] ), .Y(N326));
    AO13 un1_integ_0_0_ADD_26x26_fast_I48_Y (.A(N353), .B(integral[13])
        , .C(\un1_next_int_0_iv[13] ), .Y(N416));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I195_un1_Y (.A(N536), .B(
        \state_RNIJL492[0]_net_1 ), .Y(I195_un1_Y));
    NOR3B \state_RNI73LO3[0]  (.A(sr_new_1_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[12] ), .Y(\un2_next_int_m[12] ));
    DFN1E0C0 \integ[3]  (.D(\un1_integ[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_done), .Q(\integ[3]_net_1 ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I252_Y (.A(I174_un1_Y), .B(
        ADD_26x26_fast_I207_Y_2), .C(ADD_26x26_fast_I252_Y_0), .Y(
        \un1_integ[22] ));
    XA1A \state_RNI2U2S2[1]  (.A(sr_old_0_0), .B(\inf_abs1[3]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[3] ));
    DFN1E0C0 \integ[6]  (.D(\un1_integ[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_done), .Q(integral[6]));
    XNOR2 inf_abs0_a_0_I_14 (.A(sr_new[5]), .B(N_9_0), .Y(
        \inf_abs0_a_0[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_1 (.A(N529), .B(N514), .C(
        ADD_26x26_fast_I210_Y_0), .Y(ADD_26x26_fast_I210_Y_1));
    AND3 inf_abs0_a_0_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[5] ), .Y(
        \DWACT_FINC_E[6] ));
    NOR2 \state_RNIFJ4_0[0]  (.A(\state[1]_net_1 ), .B(
        \state[0]_net_1 ), .Y(int_done_0));
    NOR2B \state_RNI4LCR3[0]  (.A(\inf_abs0[11]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[11] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y (.A(N533), .B(I194_un1_Y), 
        .C(ADD_26x26_fast_I239_Y_0), .Y(\un1_integ[9] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_0 (.A(N399), .B(N402), .C(
        N398), .Y(ADD_26x26_fast_I206_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I58_Y (.A(N338), .B(N342), .C(
        N341), .Y(N426));
    NOR2B \state_RNILG2D[0]  (.A(sr_new[5]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[5] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I67_Y (.A(N327), .B(N330), .Y(
        N435));
    XA1A \state_RNIOF1M5[1]  (.A(sr_old[12]), .B(\inf_abs1[9]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[9] ));
    OR3 \state_RNI8RNR6[0]  (.A(\inf_abs0_m[3] ), .B(
        \un1_next_int_iv_0[3] ), .C(\un2_next_int_m[3] ), .Y(
        \un1_next_int[3] ));
    XNOR2 inf_abs0_a_0_I_12 (.A(sr_new[4]), .B(N_10), .Y(
        \inf_abs0_a_0[4] ));
    NOR2B \state_RNIV51E[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), .Y(
        next_int_0_sqmuxa_1));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I253_Y_0 (.A(integral[23]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I253_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I64_Y (.A(N329), .B(N333), .C(
        N332), .Y(N432));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I50_un1_Y (.A(N350), .B(N354), 
        .Y(I50_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I204_un1_Y_0 (.A(N502), .B(N518)
        , .Y(ADD_26x26_fast_I204_un1_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I212_un1_Y (.A(
        ADD_26x26_fast_I212_un1_Y_0), .B(N518), .Y(I212_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I127_Y (.A(N401), .B(
        ADD_26x26_fast_I127_Y_0), .C(N458), .Y(N504));
    AO1 un1_integ_0_0_ADD_26x26_fast_I110_Y (.A(N432), .B(N429), .C(
        N428), .Y(N481));
    OR2 un1_integ_0_0_ADD_26x26_fast_I90_Y (.A(N408), .B(I90_un1_Y), 
        .Y(N461));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I233_Y (.A(\un1_next_int[3] ), 
        .B(\integ[3]_net_1 ), .C(N491), .Y(\un1_integ[3] ));
    NOR3A inf_abs0_a_0_I_31 (.A(\DWACT_FINC_E[6] ), .B(sr_new[9]), .C(
        sr_new[10]), .Y(N_3_1));
    AO1B un1_integ_0_0_ADD_26x26_fast_I47_Y (.A(integral[13]), .B(
        integral[14]), .C(\un1_next_int_0_iv[13] ), .Y(N415));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I119_Y (.A(N441), .B(N437), .Y(
        N490));
    MX2 \inf_abs0[7]  (.A(sr_new[7]), .B(\inf_abs0_a_0[7] ), .S(
        sr_new_1_0), .Y(\inf_abs0[7]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I70_Y (.A(N320), .B(N324), .C(
        N323), .Y(N438));
    DFN1E0C0 \integ[5]  (.D(\un1_integ[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_done), .Q(\integ[5]_net_1 ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I44_Y (.A(integral[14]), .B(
        integral[15]), .C(\un1_next_int_0_iv_0[13] ), .Y(I90_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I245_Y (.A(N521), .B(I188_un1_Y), 
        .C(ADD_26x26_fast_I245_Y_0), .Y(\un1_integ[15] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I95_Y (.A(N413), .B(N417), .Y(
        N466));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I239_Y_0 (.A(integral[9]), .B(
        \state_RNISE23D[0]_net_1 ), .Y(ADD_26x26_fast_I239_Y_0));
    DFN1E0C0 \integ[2]  (.D(\un1_integ[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_done), .Q(\integ[2]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I135_Y (.A(N466), .B(N458), .Y(
        N512));
    OR2 un1_integ_0_0_ADD_26x26_fast_I88_Y (.A(N410), .B(N406), .Y(
        N459));
    AX1D un1_integ_0_0_ADD_26x26_fast_I247_Y (.A(I212_un1_Y), .B(
        ADD_26x26_fast_I212_Y_0), .C(ADD_26x26_fast_I247_Y_0), .Y(
        \un1_integ[17] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I237_Y_0 (.A(integral[7]), .B(
        \state_RNIU2U5B[0]_net_1 ), .Y(ADD_26x26_fast_I237_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I143_Y (.A(N466), .B(N474), .Y(
        N520));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I57_Y (.A(N345), .B(N342), .Y(
        N425));
    NOR3 inf_abs0_a_0_I_29 (.A(sr_new[7]), .B(sr_new[6]), .C(sr_new[8])
        , .Y(\DWACT_FINC_E_0[5] ));
    DFN1E0C0 \integ[23]  (.D(\un1_integ[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[23]));
    OR2 un1_integ_0_0_ADD_26x26_fast_I8_P0N (.A(integral[8]), .B(
        \un1_next_int[8] ), .Y(N342));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_2 (.A(
        ADD_26x26_fast_I206_un1_Y_0), .B(N522), .C(
        ADD_26x26_fast_I206_Y_1), .Y(ADD_26x26_fast_I206_Y_2));
    OR3 \state_RNI00AMD[0]  (.A(\inf_abs0_m[10] ), .B(
        \un1_next_int_iv_0[10] ), .C(\un2_next_int_m[10] ), .Y(
        \state_RNI00AMD[0]_net_1 ));
    INV \integ_RNIK276[25]  (.A(integral[25]), .Y(integral_i[25]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I54_Y (.A(N344), .B(N348), .C(
        N347), .Y(N422));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I131_Y (.A(N405), .B(N401), .C(
        N462), .Y(N508));
    XNOR2 inf_abs0_a_0_I_26 (.A(sr_new[9]), .B(N_5), .Y(
        \inf_abs0_a_0[9] ));
    NOR3B inf_abs1_a_1_I_19 (.A(\DWACT_FINC_E[2] ), .B(
        \DWACT_FINC_E_0[0] ), .C(sr_old[6]), .Y(N_7));
    NOR3C \state_RNIIS3M[1]  (.A(sr_old[0]), .B(\state[1]_net_1 ), .C(
        sr_old_0_0), .Y(\inf_abs1_m[0] ));
    NOR3B inf_abs1_a_1_I_16 (.A(\DWACT_FINC_E[1] ), .B(
        \DWACT_FINC_E_0[0] ), .C(sr_old[5]), .Y(N_8));
    NOR3B \state_RNIMBJV3[0]  (.A(sr_new_1_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[10]_net_1 ), .Y(\un2_next_int_m[10] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I254_Y (.A(I205_un1_Y), .B(
        ADD_26x26_fast_I205_Y_3), .C(ADD_26x26_fast_I254_Y_0), .Y(
        \un1_integ[24] ));
    DFN1E0C0 \integ[19]  (.D(\un1_integ[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[19]));
    OR3 \state_RNIJ1O9E[0]  (.A(\inf_abs0_m[11] ), .B(
        \un1_next_int_iv_0[11] ), .C(\un2_next_int_m[11] ), .Y(
        \state_RNIJ1O9E[0]_net_1 ));
    NOR2 inf_abs0_a_0_I_15 (.A(sr_new[4]), .B(sr_new[3]), .Y(
        \DWACT_FINC_E_0[1] ));
    NOR3A \state_RNIJT3M[1]  (.A(\state[1]_net_1 ), .B(sr_old_0_0), .C(
        sr_old[1]), .Y(\un18_next_int_m[1] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I161_un1_Y (.A(N486), .B(N493), 
        .Y(I161_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I117_Y (.A(N439), .B(N435), .Y(
        N488));
    OR2 \state_RNI57GE8[0]  (.A(\un1_next_int_iv_1[8] ), .B(
        \un2_next_int_m[8] ), .Y(\un1_next_int[8] ));
    DFN1E0C0 \integ[17]  (.D(\un1_integ[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[17]));
    XOR2 inf_abs0_a_0_I_5 (.A(sr_new[0]), .B(sr_new[1]), .Y(
        \inf_abs0_a_0[1] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I33_Y (.A(integral[20]), .B(
        integral[21]), .C(\un1_next_int_0_iv_0[13] ), .Y(N401));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I255_Y_0 (.A(integral[25]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I255_Y_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I127_Y_0 (.A(integral[23]), .B(
        integral[22]), .C(\un1_next_int_0_iv_0[13] ), .Y(
        ADD_26x26_fast_I127_Y_0));
    DFN1E0C0 \integ[14]  (.D(\un1_integ[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[14]));
    XNOR2 inf_abs0_a_0_I_17 (.A(sr_new[6]), .B(N_8_0), .Y(
        \inf_abs0_a_0[6] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I87_Y (.A(N405), .B(N409), .Y(
        N458));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y_0 (.A(\integ[2]_net_1 ), 
        .B(\un1_next_int[2] ), .Y(ADD_26x26_fast_I232_Y_0));
    XA1A \state_RNIB23A3[1]  (.A(sr_old_0_0), .B(\inf_abs1[4]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[4] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I84_Y (.A(N406), .B(N402), .Y(
        N455));
    AO1 un1_integ_0_0_ADD_26x26_fast_I154_Y (.A(N485), .B(N478), .C(
        N477), .Y(N531));
    MX2 \inf_abs1[11]  (.A(sr_old[11]), .B(\inf_abs1_a_1[11] ), .S(
        sr_old_0_0), .Y(\inf_abs1[11]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I11_G0N (.A(integral[11]), .B(
        \state_RNIJ1O9E[0]_net_1 ), .Y(N350));
    MX2 \inf_abs1[2]  (.A(sr_old[2]), .B(\inf_abs1_a_1[2] ), .S(
        sr_old[12]), .Y(\inf_abs1[2]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I140_Y (.A(N471), .B(N464), .C(
        N463), .Y(N517));
    OR3 \state_RNII2854[1]  (.A(\inf_abs0_m[5] ), .B(
        \un18_next_int_m[5] ), .C(\inf_abs1_m[5] ), .Y(
        \un1_next_int_iv_1[5] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I149_Y (.A(N480), .B(N472), .Y(
        N526));
    OR2 un1_integ_0_0_ADD_26x26_fast_I158_Y (.A(I158_un1_Y), .B(N481), 
        .Y(N535));
    MX2 \inf_abs1[9]  (.A(sr_old[9]), .B(\inf_abs1_a_1[9] ), .S(
        sr_old[12]), .Y(\inf_abs1[9]_net_1 ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I249_Y_0 (.A(integral[19]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I249_Y_0));
    DFN1E0C0 \integ[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done), .Q(integral[25]));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I247_Y_0 (.A(integral[17]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I247_Y_0));
    NOR3B \state_RNIJEQV1[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[3]_net_1 ), .Y(\un2_next_int_m[3] ));
    MX2 \inf_abs1[6]  (.A(sr_old[6]), .B(\inf_abs1_a_1[6] ), .S(
        sr_old[12]), .Y(\inf_abs1[6]_net_1 ));
    NOR3 inf_abs0_a_0_I_33 (.A(sr_new[10]), .B(sr_new[9]), .C(
        sr_new[11]), .Y(\DWACT_FINC_E[7] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y_0 (.A(\integ[0]_net_1 ), 
        .B(N_3), .Y(ADD_26x26_fast_I230_Y_0));
    NOR2B \state_RNI732C4[1]  (.A(\inf_abs1_a_1[8] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[8] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I242_Y (.A(N527), .B(I191_un1_Y), 
        .C(ADD_26x26_fast_I242_Y_0), .Y(\un1_integ[12] ));
    XNOR2 inf_abs0_a_0_I_20 (.A(sr_new[7]), .B(N_7_0), .Y(
        \inf_abs0_a_0[7] ));
    DFN1E0C0 \integ[11]  (.D(\un1_integ[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[11]));
    DFN1E0C0 \integ[16]  (.D(\un1_integ[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[16]));
    XNOR2 inf_abs1_a_1_I_28 (.A(sr_old[10]), .B(N_4), .Y(
        \inf_abs1_a_1[10] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_1 (.A(N516), .B(N531), .C(
        ADD_26x26_fast_I211_Y_0), .Y(ADD_26x26_fast_I211_Y_1));
    NOR3 inf_abs1_a_1_I_10 (.A(sr_old[1]), .B(sr_old[0]), .C(sr_old[2])
        , .Y(\DWACT_FINC_E_0[0] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I254_Y_0 (.A(integral[24]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I254_Y_0));
    MX2B un1_next_int_0_sqmuxa_0__m2 (.A(sr_new_0_0), .B(sr_old_0_0), 
        .S(\state[1]_net_1 ), .Y(N_3));
    OR2 un1_integ_0_0_ADD_26x26_fast_I96_Y (.A(I96_un1_Y), .B(N414), 
        .Y(N467));
    MX2 \inf_abs0[10]  (.A(sr_new[10]), .B(\inf_abs0_a_0[10] ), .S(
        sr_new_1_0), .Y(\inf_abs0[10]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I2_G0N (.A(\un1_next_int[2] ), 
        .B(\integ[2]_net_1 ), .Y(N323));
    AO1 un1_integ_0_0_ADD_26x26_fast_I114_Y (.A(N436), .B(N433), .C(
        N432), .Y(N485));
    OA1 un1_integ_0_0_ADD_26x26_fast_I189_un1_Y (.A(N485), .B(
        I161_un1_Y), .C(N524), .Y(I189_un1_Y));
    NOR2 inf_abs0_a_0_I_21 (.A(sr_new[6]), .B(sr_new[7]), .Y(
        \DWACT_FINC_E_0[3] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I147_Y (.A(N478), .B(N470), .Y(
        N524));
    DFN1E0C0 \integ[9]  (.D(\un1_integ[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_done), .Q(integral[9]));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I242_Y_0 (.A(integral[12]), .B(
        \un1_next_int[12] ), .Y(ADD_26x26_fast_I242_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I235_Y (.A(N487), .B(I162_un1_Y), 
        .C(ADD_26x26_fast_I235_Y_0), .Y(\un1_integ[5] ));
    NOR2B \state_RNIHC2D[0]  (.A(sr_new[1]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[1] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I212_Y_0 (.A(N533), .B(N518), .C(
        N517), .Y(ADD_26x26_fast_I212_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I63_Y (.A(N333), .B(N336), .Y(
        N431));
    NOR2A inf_abs1_a_1_I_11 (.A(\DWACT_FINC_E_0[0] ), .B(sr_old[3]), 
        .Y(N_10_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I96_un1_Y (.A(N418), .B(N415), 
        .Y(I96_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I118_Y (.A(I118_un1_Y), .B(N436), 
        .Y(N489));
    NOR3B \state_RNIP6T83[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[7]_net_1 ), .Y(\un2_next_int_m[7] ));
    NOR3B \state_RNI6FKU2[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[6]_net_1 ), .Y(\un2_next_int_m[6] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I237_Y (.A(N483), .B(I160_un1_Y), 
        .C(ADD_26x26_fast_I237_Y_0), .Y(\un1_integ[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I133_Y (.A(N456), .B(N464), .Y(
        N510));
    MX2 \inf_abs0[2]  (.A(sr_new[2]), .B(\inf_abs0_a_0[2] ), .S(
        sr_new_1_0), .Y(\inf_abs0[2]_net_1 ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I30_Y (.A(integral[22]), .B(
        integral[21]), .C(\un1_next_int_0_iv_0[13] ), .Y(N398));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I160_un1_Y (.A(N484), .B(N491), 
        .Y(I160_un1_Y));
    DFN1E0C0 \integ[22]  (.D(\un1_integ[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[22]));
    NOR3 inf_abs1_a_1_I_8 (.A(sr_old[1]), .B(sr_old[0]), .C(sr_old[2]), 
        .Y(N_11));
    AO1B un1_integ_0_0_ADD_26x26_fast_I43_Y (.A(integral[15]), .B(
        integral[16]), .C(\un1_next_int_0_iv_0[13] ), .Y(N411));
    NOR2 \state_RNIFJ4[0]  (.A(\state[1]_net_1 ), .B(\state[0]_net_1 ), 
        .Y(int_done));
    DFN1E0C0 \integ_0[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done), .Q(integral_0_0));
    DFN1E0C0 \integ[1]  (.D(\un1_integ[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_done), .Q(\integ[1]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I35_Y (.A(integral[20]), .B(
        integral[19]), .C(\un1_next_int_0_iv_0[13] ), .Y(N403));
    NOR2B inf_abs0_a_0_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I53_Y (.A(N348), .B(N351), .Y(
        N421));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I91_Y (.A(N413), .B(N409), .Y(
        N462));
    AX1D un1_integ_0_0_ADD_26x26_fast_I250_Y (.A(I178_un1_Y), .B(
        ADD_26x26_fast_I209_Y_1), .C(ADD_26x26_fast_I250_Y_0), .Y(
        \un1_integ[20] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I240_Y_0 (.A(integral[10]), .B(
        \state_RNI00AMD[0]_net_1 ), .Y(ADD_26x26_fast_I240_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I210_Y_0 (.A(N459), .B(I136_un1_Y)
        , .Y(ADD_26x26_fast_I210_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I71_Y (.A(N324), .B(N321), .Y(
        N439));
    DFN1E0C0 \integ[20]  (.D(\un1_integ[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[20]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I244_Y (.A(N523), .B(I189_un1_Y), 
        .C(ADD_26x26_fast_I244_Y_0), .Y(\un1_integ[14] ));
    NOR3 inf_abs1_a_1_I_29 (.A(sr_old[7]), .B(sr_old[6]), .C(sr_old[8])
        , .Y(\DWACT_FINC_E[5] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I207_Y_1 (.A(N404), .B(N400), .C(
        N461), .Y(ADD_26x26_fast_I207_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I106_Y (.A(N428), .B(N425), .C(
        N424), .Y(N477));
    XNOR2 inf_abs0_a_0_I_32 (.A(sr_new[11]), .B(N_3_1), .Y(
        \inf_abs0_a_0[11] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_1 (.A(
        ADD_26x26_fast_I208_un1_Y_0), .B(N526), .C(
        ADD_26x26_fast_I208_Y_0), .Y(ADD_26x26_fast_I208_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I102_Y (.A(N424), .B(N421), .C(
        N420), .Y(N473));
    AX1D un1_integ_0_0_ADD_26x26_fast_I251_Y (.A(I176_un1_Y), .B(
        ADD_26x26_fast_I208_Y_1), .C(ADD_26x26_fast_I251_Y_0), .Y(
        \un1_integ[21] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I121_un1_Y (.A(N441), .B(
        \state_RNIJL492[0]_net_1 ), .Y(I121_un1_Y));
    XNOR2 inf_abs1_a_1_I_26 (.A(sr_old[9]), .B(N_5_0), .Y(
        \inf_abs1_a_1[9] ));
    DFN1E0C0 \integ[18]  (.D(\un1_integ[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_done_0), .Q(integral[18]));
    OR2 un1_integ_0_0_ADD_26x26_fast_I4_P0N (.A(\integ[4]_net_1 ), .B(
        \un1_next_int[4] ), .Y(N330));
    AO1 un1_integ_0_0_ADD_26x26_fast_I144_Y (.A(N475), .B(N468), .C(
        N467), .Y(N521));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I139_Y (.A(N470), .B(N462), .Y(
        N516));
    OR3 \state_RNINUFN2[0]  (.A(\un18_next_int_m[1] ), .B(
        \inf_abs1_m[1] ), .C(\un2_next_int_m[1] ), .Y(
        \un1_next_int_iv_1[1] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_0 (.A(N465), .B(N458), .C(
        N457), .Y(ADD_26x26_fast_I209_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I148_Y (.A(I148_un1_Y), .B(N471), 
        .Y(N525));
    XA1A \state_RNI0E364[1]  (.A(sr_old_0_0), .B(\inf_abs1[6]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[6] ));
    NOR2B \state_RNI6FKU2_0[0]  (.A(\inf_abs0[6]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[6] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I60_Y (.A(N335), .B(N339), .C(
        N338), .Y(N428));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y (.A(
        ADD_26x26_fast_I232_Y_0), .B(N493), .Y(\un1_integ[2] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I204_Y_2 (.A(N398), .B(
        ADD_26x26_fast_I204_Y_0), .C(N455), .Y(ADD_26x26_fast_I204_Y_2)
        );
    DFN1C0 \state[1]  (.D(\state_RNO_4[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[1]_net_1 ));
    XNOR2 inf_abs0_a_0_I_23 (.A(sr_new[8]), .B(N_6_0), .Y(
        \inf_abs0_a_0[8] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I118_un1_Y (.A(N440), .B(N437), 
        .Y(I118_un1_Y));
    NOR3A inf_abs1_a_1_I_13 (.A(\DWACT_FINC_E_0[0] ), .B(sr_old[3]), 
        .C(sr_old[4]), .Y(N_9));
    MX2 \inf_abs1[7]  (.A(sr_old[7]), .B(\inf_abs1_a_1[7] ), .S(
        sr_old[12]), .Y(\inf_abs1[7]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I9_G0N (.A(integral[9]), .B(
        \state_RNISE23D[0]_net_1 ), .Y(N344));
    OA1B un1_integ_0_0_ADD_26x26_fast_I40_Y (.A(integral[17]), .B(
        integral[16]), .C(\un1_next_int_0_iv_0[13] ), .Y(N408));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I65_Y (.A(N330), .B(N333), .Y(
        N433));
    OA1 un1_integ_0_0_ADD_26x26_fast_I207_un1_Y_0 (.A(N485), .B(
        I161_un1_Y), .C(N508), .Y(ADD_26x26_fast_I207_un1_Y_0));
    NOR3 inf_abs0_a_0_I_8 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2]), 
        .Y(N_11_0));
    AND3 inf_abs1_a_1_I_30 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E_0[6] ));
    MX2 \inf_abs1[3]  (.A(sr_old[3]), .B(\inf_abs1_a_1[3] ), .S(
        sr_old[12]), .Y(\inf_abs1[3]_net_1 ));
    XNOR2 inf_abs0_a_0_I_35 (.A(sr_new[12]), .B(N_2), .Y(
        \inf_abs0_a_0[12] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I178_un1_Y (.A(N527), .B(N512), 
        .Y(I178_un1_Y));
    OR2 \state_RNITUJS9[0]  (.A(\un1_next_int_iv_0[12] ), .B(
        \un2_next_int_m[12] ), .Y(\un1_next_int[12] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I45_Y (.A(integral[14]), .B(
        integral[15]), .C(\un1_next_int_0_iv[13] ), .Y(N413));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I137_Y (.A(N468), .B(N460), .Y(
        N514));
    OR2 \state_RNISE23D[0]  (.A(\un1_next_int_iv_1[9] ), .B(
        \un2_next_int_m[9] ), .Y(\state_RNISE23D[0]_net_1 ));
    XNOR2 inf_abs0_a_0_I_9 (.A(sr_new[3]), .B(N_11_0), .Y(
        \inf_abs0_a_0[3] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I3_P0N (.A(\integ[3]_net_1 ), .B(
        \un1_next_int[3] ), .Y(N327));
    NOR2B \state_RNO[0]  (.A(calc_int), .B(int_done), .Y(
        \state_RNO_3[0] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I50_Y (.A(I50_un1_Y), .B(N353), 
        .Y(N418));
    AO1 un1_integ_0_0_ADD_26x26_fast_I204_Y_3 (.A(N517), .B(N502), .C(
        ADD_26x26_fast_I204_Y_2), .Y(ADD_26x26_fast_I204_Y_3));
    XNOR2 inf_abs1_a_1_I_20 (.A(sr_old[7]), .B(N_7), .Y(
        \inf_abs1_a_1[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I74_un1_Y (.A(N318), .B(
        \state_RNIJL492[0]_net_1 ), .Y(I74_un1_Y));
    NOR3B \state_RNIGB2D[0]  (.A(\state[0]_net_1 ), .B(sr_new[12]), .C(
        sr_new[0]), .Y(\un2_next_int_m[0] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I36_Y (.A(integral[19]), .B(
        integral[18]), .C(\un1_next_int_0_iv_0[13] ), .Y(N404));
    NOR3A inf_abs1_a_1_I_31 (.A(\DWACT_FINC_E_0[6] ), .B(sr_old[9]), 
        .C(sr_old[10]), .Y(N_3_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I136_un1_Y (.A(N467), .B(N460), 
        .Y(I136_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I0_P0N (.A(\integ[0]_net_1 ), .B(
        N_3), .Y(N318));
    NOR2 inf_abs1_a_1_I_6 (.A(sr_old[0]), .B(sr_old[1]), .Y(N_12_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I55_Y (.A(N345), .B(N348), .Y(
        N423));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I205_un1_Y (.A(N520), .B(N504), 
        .C(N658), .Y(I205_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I163_un1_Y (.A(N490), .B(
        \state_RNIJL492[0]_net_1 ), .Y(I163_un1_Y));
    NOR2B \state_RNIJEQV1_0[0]  (.A(next_int_1_sqmuxa), .B(
        \inf_abs0[3]_net_1 ), .Y(\inf_abs0_m[3] ));
    NOR2 inf_abs1_a_1_I_21 (.A(sr_old[6]), .B(sr_old[7]), .Y(
        \DWACT_FINC_E[3] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_1 (.A(N459), .B(N452), .C(
        ADD_26x26_fast_I206_Y_0), .Y(ADD_26x26_fast_I206_Y_1));
    OA1 un1_integ_0_0_ADD_26x26_fast_I5_G0N (.A(\un2_next_int_m[5] ), 
        .B(\un1_next_int_iv_1[5] ), .C(\integ[5]_net_1 ), .Y(N332));
    AND3 inf_abs0_a_0_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(
        \DWACT_FINC_E[4] ));
    DFN1E0C0 \integ[7]  (.D(\un1_integ[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_done), .Q(integral[7]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_2 (.A(
        ADD_26x26_fast_I207_un1_Y_0), .B(N524), .C(
        ADD_26x26_fast_I207_Y_1), .Y(ADD_26x26_fast_I207_Y_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I4_G0N (.A(\integ[4]_net_1 ), 
        .B(\un1_next_int[4] ), .Y(N329));
    OR2 \state_RNI42RG_0[1]  (.A(next_int_0_sqmuxa_1), .B(
        next_int_1_sqmuxa), .Y(\un1_next_int_0_iv[13] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I195_Y (.A(I195_un1_Y), .B(N535), 
        .Y(N658));
    OA1 un1_integ_0_0_ADD_26x26_fast_I206_un1_Y_0 (.A(N483), .B(
        I160_un1_Y), .C(N506), .Y(ADD_26x26_fast_I206_un1_Y_0));
    XNOR2 inf_abs1_a_1_I_14 (.A(sr_old[5]), .B(N_9), .Y(
        \inf_abs1_a_1[5] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I234_Y (.A(N489), .B(I163_un1_Y), 
        .C(ADD_26x26_fast_I234_Y_0), .Y(\un1_integ[4] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I205_Y_2 (.A(N400), .B(
        ADD_26x26_fast_I205_Y_0), .C(N457), .Y(ADD_26x26_fast_I205_Y_2)
        );
    NOR2B un1_integ_0_0_ADD_26x26_fast_I174_un1_Y (.A(N508), .B(N523), 
        .Y(I174_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I162_un1_Y (.A(N488), .B(N442), 
        .Y(I162_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I240_Y (.A(N531), .B(I193_un1_Y), 
        .C(ADD_26x26_fast_I240_Y_0), .Y(\un1_integ[10] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I156_Y (.A(N487), .B(N480), .C(
        N479), .Y(N533));
    NOR3B \state_RNICB7V2[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[8] ), .Y(\un2_next_int_m[8] ));
    DFN1E0C0 \integ[8]  (.D(\un1_integ[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_done), .Q(integral[8]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I85_Y (.A(N407), .B(N403), .Y(
        N456));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I251_Y_0 (.A(integral[21]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I251_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I152_Y (.A(N483), .B(N476), .C(
        N475), .Y(N529));
    AND3 inf_abs0_a_0_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(N_6_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I9_P0N (.A(integral[9]), .B(
        \state_RNISE23D[0]_net_1 ), .Y(N345));
    OA1 un1_integ_0_0_ADD_26x26_fast_I208_un1_Y_0 (.A(N487), .B(
        I162_un1_Y), .C(N510), .Y(ADD_26x26_fast_I208_un1_Y_0));
    NOR2B \state_RNIP6T83_0[0]  (.A(\inf_abs0[7]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[7] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I31_Y (.A(integral[21]), .B(
        integral[22]), .C(\un1_next_int_0_iv_0[13] ), .Y(N399));
    XNOR2 inf_abs1_a_1_I_12 (.A(sr_old[4]), .B(N_10_0), .Y(
        \inf_abs1_a_1[4] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I235_Y_0 (.A(\un2_next_int_m[5] )
        , .B(\un1_next_int_iv_1[5] ), .C(\integ[5]_net_1 ), .Y(
        ADD_26x26_fast_I235_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I241_Y (.A(N529), .B(I192_un1_Y), 
        .C(ADD_26x26_fast_I241_Y_0), .Y(\un1_integ[11] ));
    NOR3 inf_abs0_a_0_I_18 (.A(sr_new[5]), .B(sr_new[4]), .C(sr_new[3])
        , .Y(\DWACT_FINC_E_0[2] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I11_P0N (.A(integral[11]), .B(
        \state_RNIJ1O9E[0]_net_1 ), .Y(N351));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I243_Y_0 (.A(integral[13]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I243_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I105_Y (.A(N423), .B(N427), .Y(
        N476));
    AO1 un1_integ_0_0_ADD_26x26_fast_I213_Y_0 (.A(N535), .B(N520), .C(
        N519), .Y(ADD_26x26_fast_I213_Y_0));
    MX2 \inf_abs0[11]  (.A(sr_new[11]), .B(\inf_abs0_a_0[11] ), .S(
        sr_new_1_0), .Y(\inf_abs0[11]_net_1 ));
    XOR2 inf_abs1_a_1_I_5 (.A(sr_old[0]), .B(sr_old[1]), .Y(
        \inf_abs1_a_1[1] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I101_Y (.A(N423), .B(N419), .Y(
        N472));
    AO1 un1_integ_0_0_ADD_26x26_fast_I66_Y (.A(N326), .B(N330), .C(
        N329), .Y(N434));
    AX1D un1_integ_0_0_ADD_26x26_fast_I248_Y (.A(I211_un1_Y), .B(
        ADD_26x26_fast_I211_Y_1), .C(ADD_26x26_fast_I248_Y_0), .Y(
        \un1_integ[18] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I99_Y (.A(N417), .B(N421), .Y(
        N470));
    OR2 un1_integ_0_0_ADD_26x26_fast_I92_Y (.A(N410), .B(N414), .Y(
        N463));
    OA1 un1_integ_0_0_ADD_26x26_fast_I191_un1_Y (.A(N489), .B(
        I163_un1_Y), .C(N528), .Y(I191_un1_Y));
    NOR2B \state_RNI4RHL1[0]  (.A(\inf_abs0[2]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[2] ));
    XA1A \state_RNI4I1U5[1]  (.A(sr_old[12]), .B(\inf_abs1[10]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[10] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I72_Y (.A(N317), .B(N321), .C(
        N320), .Y(N440));
    OA1B un1_integ_0_0_ADD_26x26_fast_I46_Y (.A(integral[13]), .B(
        integral[14]), .C(\un1_next_int_0_iv[13] ), .Y(N414));
    NOR3B \state_RNI9DJ11[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[2] ), .Y(\un2_next_int_m[2] ));
    NOR3 inf_abs1_a_1_I_33 (.A(sr_old[10]), .B(sr_old[9]), .C(
        sr_old[11]), .Y(\DWACT_FINC_E_0[7] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I116_Y (.A(N438), .B(N435), .C(
        N434), .Y(N487));
    AO1 un1_integ_0_0_ADD_26x26_fast_I112_Y (.A(N434), .B(N431), .C(
        N430), .Y(N483));
    NOR2A inf_abs0_a_0_I_25 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .Y(
        N_5));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I8_G0N (.A(integral[8]), .B(
        \un1_next_int[8] ), .Y(N341));
    MX2 \inf_abs0[3]  (.A(sr_new[3]), .B(\inf_abs0_a_0[3] ), .S(
        sr_new_1_0), .Y(\inf_abs0[3]_net_1 ));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I210_un1_Y (.A(N514), .B(N491), 
        .C(N530), .Y(I210_un1_Y));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y_0 (.A(\integ[4]_net_1 ), 
        .B(\un1_next_int[4] ), .Y(ADD_26x26_fast_I234_Y_0));
    NOR3A inf_abs0_a_0_I_27 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .C(
        sr_new[9]), .Y(N_4_0));
    
endmodule


module error_calc_13s_12s_4_1(
       cur_error,
       LED_FB_i_0,
       LED_FB,
       average,
       calc_error,
       n_rst_c,
       clk_c
    );
output [12:0] cur_error;
input  LED_FB_i_0;
input  [7:0] LED_FB;
input  [6:2] average;
input  calc_error;
input  n_rst_c;
input  clk_c;

    wire N_40, N_38, GND, VCC;
    
    AX1B un2_diffreg_1_m37 (.A(LED_FB[5]), .B(LED_FB[6]), .C(LED_FB[7])
        , .Y(N_38));
    DFN1E1C0 \diffreg[3]  (.D(average[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[3]));
    XNOR2 un2_diffreg_1_m39 (.A(LED_FB[6]), .B(LED_FB[5]), .Y(N_40));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \diffreg[7]  (.D(LED_FB[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[7]));
    DFN1E1C0 \diffreg[1]  (.D(average[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[1]));
    DFN1E1C0 \diffreg[12]  (.D(N_38), .CLK(clk_c), .CLR(n_rst_c), .E(
        calc_error), .Q(cur_error[12]));
    DFN1E1C0 \diffreg[11]  (.D(N_40), .CLK(clk_c), .CLR(n_rst_c), .E(
        calc_error), .Q(cur_error[11]));
    GND GND_i (.Y(GND));
    DFN1E1C0 \diffreg[9]  (.D(LED_FB[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[9]));
    DFN1E1C0 \diffreg[8]  (.D(LED_FB[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[8]));
    DFN1E1C0 \diffreg[6]  (.D(LED_FB[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[6]));
    DFN1E1C0 \diffreg[10]  (.D(LED_FB_i_0), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[10]));
    DFN1E1C0 \diffreg[5]  (.D(LED_FB[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[5]));
    DFN1E1C0 \diffreg[4]  (.D(average[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[4]));
    DFN1E1C0 \diffreg[2]  (.D(average[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[2]));
    DFN1E1C0 \diffreg[0]  (.D(average[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[0]));
    
endmodule


module derivative_calc_13s_4_1(
       derivative_0,
       sr_new,
       sr_prev,
       deriv_enable,
       n_rst_c,
       clk_c
    );
output derivative_0;
input  [12:0] sr_new;
input  [12:0] sr_prev;
input  deriv_enable;
input  n_rst_c;
input  clk_c;

    wire SUB_13x13_medium_area_I49_Y_1, N208, N176, 
        SUB_13x13_medium_area_I49_Y_0, 
        SUB_13x13_medium_area_I26_un1_Y_0, 
        SUB_13x13_medium_area_I49_un1_Y_1, 
        SUB_13x13_medium_area_I49_un1_Y_0, N_15, 
        SUB_13x13_medium_area_I42_Y_1, N218, N180, 
        SUB_13x13_medium_area_I42_Y_0, 
        SUB_13x13_medium_area_I30_un1_Y_0, 
        SUB_13x13_medium_area_I42_un1_Y_1, 
        SUB_13x13_medium_area_I42_un1_Y_0, N_7, 
        SUB_13x13_medium_area_I41_Y_0, 
        SUB_13x13_medium_area_I34_un1_Y_0, 
        SUB_13x13_medium_area_I41_un1_Y_0, N_5, 
        SUB_13x13_medium_area_I28_un1_Y_0, 
        SUB_13x13_medium_area_I32_un1_Y_0, N204, N212, N_24, N226, 
        N222, N185, N_13, N_21, GND, VCC;
    
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I34_un1_Y_0 (.A(
        sr_new[1]), .B(sr_prev[1]), .Y(
        SUB_13x13_medium_area_I34_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y_0 (.A(
        SUB_13x13_medium_area_I30_un1_Y_0), .B(sr_new[6]), .C(
        sr_prev[6]), .Y(SUB_13x13_medium_area_I42_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I15_S (.A(sr_new[2]), 
        .B(sr_prev[2]), .Y(N_5));
    OR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I36_Y (.A(sr_prev[0]), 
        .B(sr_new[0]), .Y(N185));
    XNOR3 un2_deriv_out_0_0_SUB_13x13_medium_area_I82_Y (.A(sr_new[12])
        , .B(sr_prev[12]), .C(N226), .Y(N_24));
    VCC VCC_i (.Y(VCC));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I64_Y (.A(N204), .B(
        sr_new[11]), .C(sr_prev[11]), .Y(N226));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I41_Y_0 (.A(
        SUB_13x13_medium_area_I34_un1_Y_0), .B(sr_new[2]), .C(
        sr_prev[2]), .Y(SUB_13x13_medium_area_I41_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I19_S (.A(sr_prev[6]), 
        .B(sr_new[6]), .Y(N_13));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I42_un1_Y_0 (.A(
        sr_new[4]), .B(sr_prev[4]), .C(N_7), .Y(
        SUB_13x13_medium_area_I42_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I28_Y (.A(
        SUB_13x13_medium_area_I28_un1_Y_0), .B(sr_new[8]), .C(
        sr_prev[8]), .Y(N208));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y_1 (.A(N218), .B(
        N180), .C(SUB_13x13_medium_area_I42_Y_0), .Y(
        SUB_13x13_medium_area_I42_Y_1));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I28_un1_Y_0 (.A(
        sr_new[7]), .B(sr_prev[7]), .Y(
        SUB_13x13_medium_area_I28_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y_0 (.A(
        SUB_13x13_medium_area_I26_un1_Y_0), .B(sr_new[10]), .C(
        sr_prev[10]), .Y(SUB_13x13_medium_area_I49_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I20_S (.A(sr_new[7]), 
        .B(sr_prev[7]), .Y(N_15));
    DFN1E1C0 \deriv_out[12]  (.D(N_24), .CLK(clk_c), .CLR(n_rst_c), .E(
        deriv_enable), .Q(derivative_0));
    GND GND_i (.Y(GND));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I23_S (.A(sr_new[10]), 
        .B(sr_prev[10]), .Y(N_21));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I26_un1_Y_0 (.A(
        sr_new[9]), .B(sr_prev[9]), .Y(
        SUB_13x13_medium_area_I26_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I32_Y (.A(
        SUB_13x13_medium_area_I32_un1_Y_0), .B(sr_new[4]), .C(
        sr_prev[4]), .Y(N218));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I30_un1_Y_0 (.A(
        sr_new[5]), .B(sr_prev[5]), .Y(
        SUB_13x13_medium_area_I30_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y (.A(
        SUB_13x13_medium_area_I49_un1_Y_1), .B(N212), .C(
        SUB_13x13_medium_area_I49_Y_1), .Y(N204));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I32_un1_Y_0 (.A(
        sr_new[3]), .B(sr_prev[3]), .Y(
        SUB_13x13_medium_area_I32_un1_Y_0));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I31_Y (.A(sr_new[5]), 
        .B(sr_prev[5]), .C(N_13), .Y(N180));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I41_un1_Y_0 (.A(
        sr_new[1]), .B(sr_prev[1]), .C(N_5), .Y(
        SUB_13x13_medium_area_I41_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y_1 (.A(N208), .B(
        N176), .C(SUB_13x13_medium_area_I49_Y_0), .Y(
        SUB_13x13_medium_area_I49_Y_1));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I16_S (.A(sr_prev[3]), 
        .B(sr_new[3]), .Y(N_7));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y (.A(
        SUB_13x13_medium_area_I42_un1_Y_1), .B(N222), .C(
        SUB_13x13_medium_area_I42_Y_1), .Y(N212));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I27_Y (.A(sr_new[9]), 
        .B(sr_prev[9]), .C(N_21), .Y(N176));
    NOR2B un2_deriv_out_0_0_SUB_13x13_medium_area_I49_un1_Y_1 (.A(
        SUB_13x13_medium_area_I49_un1_Y_0), .B(N176), .Y(
        SUB_13x13_medium_area_I49_un1_Y_1));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I49_un1_Y_0 (.A(
        sr_prev[8]), .B(sr_new[8]), .C(N_15), .Y(
        SUB_13x13_medium_area_I49_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I41_Y (.A(
        SUB_13x13_medium_area_I41_un1_Y_0), .B(N185), .C(
        SUB_13x13_medium_area_I41_Y_0), .Y(N222));
    NOR2B un2_deriv_out_0_0_SUB_13x13_medium_area_I42_un1_Y_1 (.A(
        SUB_13x13_medium_area_I42_un1_Y_0), .B(N180), .Y(
        SUB_13x13_medium_area_I42_un1_Y_1));
    
endmodule


module pwm_tx_400s_32s_13s_10_1000000s_45s_1_0(
       off_div,
       act_ctl_5_i,
       act_ctl_5_3,
       act_ctl_5_0,
       pwm_chg_0,
       pwm_chg,
       n_rst_c,
       clk_c,
       act_ctl_5_2,
       act_ctl_5_1,
       act_ctl_5_9,
       act_ctl_5_8,
       act_ctl_5,
       primary_fb_c
    );
input  [31:0] off_div;
input  act_ctl_5_i;
input  act_ctl_5_3;
input  act_ctl_5_0;
input  pwm_chg_0;
input  pwm_chg;
input  n_rst_c;
input  clk_c;
input  act_ctl_5_2;
input  act_ctl_5_1;
input  act_ctl_5_9;
input  act_ctl_5_8;
input  act_ctl_5;
output primary_fb_c;

    wire N_400_0, I_140_4, I_140_3, \DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] , \DWACT_COMP0_E[1] , N_18, 
        I_20_4, \counter[7]_net_1 , N_20, I_23_6, \counter[8]_net_1 , 
        N_11, N_6, N_8, \DWACT_FDEC_E[0] , N_3, \DWACT_FDEC_E[2] , 
        N_16, N_14, \counter[6]_net_1 , N_2, \counter[2]_net_1 , 
        counter_m6_0_a2_7, counter_m6_0_a2_2, counter_m6_0_a2_1, 
        counter_m6_0_a2_6, \counter[16]_net_1 , \counter[18]_net_1 , 
        counter_m6_0_a2_4, \counter[15]_net_1 , \counter[10]_net_1 , 
        \counter[17]_net_1 , \counter[13]_net_1 , \counter[14]_net_1 , 
        \counter[11]_net_1 , \counter[12]_net_1 , counter_c18, 
        \counter[9]_net_1 , counter_c8, counter_n31, 
        \counter[31]_net_1 , counter_63_0, cur_pwm_RNIVKRSJ2_0_net_1, 
        \counter[30]_net_1 , counter_c29, counter_n30, counter_n29, 
        \counter[29]_net_1 , counter_c28, counter_n28, counter_n28_tz, 
        \counter[27]_net_1 , counter_c26, \counter[28]_net_1 , 
        counter_n27, counter_n26, counter_n26_tz, \counter[25]_net_1 , 
        counter_c24, \counter[26]_net_1 , counter_n25, counter_n24, 
        counter_n24_tz, \counter[23]_net_1 , counter_c22, 
        \counter[24]_net_1 , counter_n23, counter_n22, counter_n22_tz, 
        \counter[21]_net_1 , counter_c20, \counter[22]_net_1 , 
        counter_n21, counter_n20, counter_n20_tz, \counter[19]_net_1 , 
        \counter[20]_net_1 , counter_n19, counter_n18, counter_c17, 
        counter_n17, counter_c16, counter_n16, counter_c15, 
        counter_n15, counter_c14, counter_n14, counter_c13, 
        counter_n13, counter_c12, counter_n12, counter_c11, 
        counter_n11, counter_c10, counter_n10, counter_n10_tz, 
        counter_n9, counter_n8, counter_n8_tz, counter_c6, counter_n7, 
        counter_n6, counter_n6_tz, \counter[5]_net_1 , counter_c4, 
        counter_n5, counter_n4, counter_n4_tz, \counter[3]_net_1 , 
        counter_c2, \counter[4]_net_1 , counter_n3, counter_n2, 
        counter_n2_tz, \counter[1]_net_1 , \counter[0]_net_1 , 
        \off_time[0] , \off_reg[0]_net_1 , \off_time[1] , 
        \off_reg[1]_net_1 , \off_time[3] , \off_reg[3]_net_1 , 
        \off_time[4] , \off_reg[4]_net_1 , \off_time[8] , 
        \off_reg[8]_net_1 , \off_time[10] , \off_reg[10]_net_1 , 
        \off_time[11] , \off_reg[11]_net_1 , \off_time[12] , 
        \off_reg[12]_net_1 , \off_time[17] , \off_reg[17]_net_1 , 
        \off_time[20] , \off_reg[20]_net_1 , \off_time[23] , 
        \off_reg[23]_net_1 , \off_time[18] , \off_reg[18]_net_1 , 
        \off_time[26] , \off_reg[26]_net_1 , \off_time[9] , 
        \off_reg[9]_net_1 , \off_time[21] , \off_reg[21]_net_1 , 
        \off_time[5] , \off_reg[5]_net_1 , \off_time[14] , 
        \off_reg[14]_net_1 , \off_time[16] , \off_reg[16]_net_1 , 
        \off_time[25] , \off_reg[25]_net_1 , \off_time[22] , 
        \off_reg[22]_net_1 , \off_time[27] , \off_reg[27]_net_1 , 
        \off_time[31] , \off_reg[31]_net_1 , \off_time[29] , 
        \off_reg[29]_net_1 , \off_time[30] , \off_reg[30]_net_1 , 
        \off_time[28] , \off_reg[28]_net_1 , \off_time[24] , 
        \off_reg[24]_net_1 , \off_time[15] , \off_reg[15]_net_1 , 
        \off_time[13] , \off_reg[13]_net_1 , \off_time[7] , 
        \off_reg[7]_net_1 , \off_time[6] , \off_reg[6]_net_1 , 
        \off_time[19] , \off_reg[19]_net_1 , \off_time[2] , 
        \off_reg[2]_net_1 , counter_n1, \counter_RNO_1[0] , 
        cur_pwm_RNO_1, \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] , N_4, N_21, N_17, N_13, 
        I_14_4, \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] , \DWACT_BL_EQUAL_0_E[3] , 
        \DWACT_BL_EQUAL_0_E[2] , \DWACT_BL_EQUAL_0_E[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] , \DWACT_COMP0_E_0[1] , 
        \DWACT_COMP0_E_0[2] , \DWACT_COMP0_E[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] , N_11_0, N_10, N_9, N_6_0, 
        N_8_0, N_7, N_5, N_2_0, N_3_0, N_4_0, N_21_0, N_20_0, N_19, 
        N_16_0, N_18_0, N_17_0, N_15, N_12, N_13_0, N_14_0, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] , 
        \DWACT_BL_EQUAL_0_E[4] , \DWACT_BL_EQUAL_0_E_0[3] , 
        \DWACT_BL_EQUAL_0_E_0[0] , \DWACT_BL_EQUAL_0_E[1] , 
        \DWACT_BL_EQUAL_0_E_0[2] , \DWACT_CMPLE_PO0_DWACT_COMP0_E[1] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[0] , N_31, N_30, N_29, N_26, 
        N_28, N_27, N_25, N_22, N_23, N_24, \ACT_LT4_E[3] , 
        \ACT_LT4_E[6] , \ACT_LT4_E[10] , \ACT_LT4_E[7] , 
        \ACT_LT4_E[8] , \ACT_LT4_E[5] , \ACT_LT4_E[4] , \ACT_LT4_E[0] , 
        \ACT_LT4_E[1] , \ACT_LT4_E[2] , \DWACT_BL_EQUAL_0_E_1[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] , 
        \DWACT_BL_EQUAL_0_E_1[0] , \DWACT_BL_EQUAL_0_E_0[1] , 
        \DWACT_BL_EQUAL_0_E_1[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] , 
        \DWACT_BL_EQUAL_0_E_2[0] , \DWACT_BL_EQUAL_0_E_1[1] , 
        \DWACT_BL_EQUAL_0_E_2[2] , \DWACT_BL_EQUAL_0_E_2[3] , 
        \DWACT_BL_EQUAL_0_E_0[4] , \DWACT_BL_EQUAL_0_E[5] , 
        \DWACT_BL_EQUAL_0_E[6] , \DWACT_BL_EQUAL_0_E[7] , 
        \DWACT_BL_EQUAL_0_E[8] , \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] , N_41, N_40, N_39, N_36, 
        N_38, N_37, N_35, N_32, N_33, N_34, \ACT_LT3_E[3] , 
        \ACT_LT3_E[4] , \ACT_LT3_E[5] , \ACT_LT3_E[0] , \ACT_LT3_E[1] , 
        \ACT_LT3_E[2] , \DWACT_BL_EQUAL_0_E_3[2] , 
        \DWACT_BL_EQUAL_0_E_2[1] , \DWACT_BL_EQUAL_0_E_3[0] , N_51, 
        N_50, N_49, N_46, N_48, N_47, N_45, N_42, N_43, N_44, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] , 
        \DWACT_BL_EQUAL_0_E_1[4] , \DWACT_BL_EQUAL_0_E_3[3] , 
        \DWACT_BL_EQUAL_0_E_4[0] , \DWACT_BL_EQUAL_0_E_3[1] , 
        \DWACT_BL_EQUAL_0_E_4[2] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] , 
        \DWACT_BL_EQUAL_0_E[12] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] , 
        \DWACT_BL_EQUAL_0_E_5[0] , \DWACT_BL_EQUAL_0_E_4[1] , 
        \DWACT_BL_EQUAL_0_E_5[2] , \DWACT_BL_EQUAL_0_E_4[3] , 
        \DWACT_BL_EQUAL_0_E_2[4] , \DWACT_BL_EQUAL_0_E_0[5] , 
        \DWACT_BL_EQUAL_0_E_0[6] , \DWACT_BL_EQUAL_0_E_0[7] , 
        \DWACT_BL_EQUAL_0_E_0[8] , \DWACT_BL_EQUAL_0_E[9] , 
        \DWACT_BL_EQUAL_0_E[10] , \DWACT_BL_EQUAL_0_E[11] , N_2_1, 
        N_5_0, GND, VCC;
    
    DFN1C0 \counter[19]  (.D(counter_n19), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[19]_net_1 ));
    AND3 un1_counter_0_I_78 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] ));
    NOR3 un1_counter_2_0_I_17 (.A(\counter[20]_net_1 ), .B(
        \counter[19]_net_1 ), .C(\counter[21]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] ));
    XOR2 un1_act_ctl_I_23 (.A(act_ctl_5), .B(N_2_1), .Y(I_23_6));
    NOR2A \off_reg_RNIQ089[27]  (.A(\off_reg[27]_net_1 ), .B(
        act_ctl_5_2), .Y(\off_time[27] ));
    AND2A un1_counter_0_I_51 (.A(\off_time[26] ), .B(
        \counter[26]_net_1 ), .Y(\ACT_LT3_E[5] ));
    NOR3C \counter_RNI9EN95[19]  (.A(\counter[19]_net_1 ), .B(
        counter_c18), .C(\counter[20]_net_1 ), .Y(counter_c20));
    NOR2A \off_reg_RNIDSPM[5]  (.A(\off_reg[5]_net_1 ), .B(act_ctl_5_9)
        , .Y(\off_time[5] ));
    DFN1E1C0 \off_reg[28]  (.D(off_div[28]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[28]_net_1 ));
    AX1C \counter_RNO_0[2]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .C(\counter[2]_net_1 ), .Y(counter_n2_tz));
    DFN1C0 \counter[28]  (.D(counter_n28), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[28]_net_1 ));
    XNOR2 un1_counter_0_I_73 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .Y(\DWACT_BL_EQUAL_0_E_2[2] ));
    OA1A un1_counter_0_I_136 (.A(N_6_0), .B(N_8_0), .C(N_7), .Y(N_11_0)
        );
    NOR2A \off_reg_RNIS289[29]  (.A(\off_reg[29]_net_1 ), .B(
        act_ctl_5_2), .Y(\off_time[29] ));
    OA1A un1_counter_0_I_132 (.A(\counter[3]_net_1 ), .B(\off_time[3] )
        , .C(N_3_0), .Y(N_7));
    DFN1E1C0 \off_reg[15]  (.D(off_div[15]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[15]_net_1 ));
    DFN1E1C0 \off_reg[26]  (.D(off_div[26]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[26]_net_1 ));
    AND3 un1_counter_0_I_14 (.A(\DWACT_BL_EQUAL_0_E[9] ), .B(
        \DWACT_BL_EQUAL_0_E[10] ), .C(\DWACT_BL_EQUAL_0_E[11] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] ));
    NOR2A \off_reg_RNI9MML[2]  (.A(\off_reg[2]_net_1 ), .B(act_ctl_5_8)
        , .Y(\off_time[2] ));
    XA1B \counter_RNO[11]  (.A(\counter[11]_net_1 ), .B(counter_c10), 
        .C(N_400_0), .Y(counter_n11));
    DFN1C0 \counter[29]  (.D(counter_n29), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[29]_net_1 ));
    DFN1E1C0 \off_reg[5]  (.D(off_div[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[5]_net_1 ));
    NOR3 un1_counter_2_0_I_77 (.A(\counter[12]_net_1 ), .B(
        \counter[10]_net_1 ), .C(\counter[11]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] ));
    XNOR2 un1_counter_0_I_82 (.A(\counter[15]_net_1 ), .B(
        \off_time[15] ), .Y(\DWACT_BL_EQUAL_0_E_1[0] ));
    DFN1C0 \counter[11]  (.D(counter_n11), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[11]_net_1 ));
    XNOR2 un1_counter_0_I_109 (.A(\counter[6]_net_1 ), .B(
        \off_time[6] ), .Y(\DWACT_BL_EQUAL_0_E[1] ));
    NOR2A \off_reg_RNIMP38[15]  (.A(\off_reg[15]_net_1 ), .B(
        act_ctl_5_1), .Y(\off_time[15] ));
    NOR2A \off_reg_RNI8LML[1]  (.A(\off_reg[1]_net_1 ), .B(act_ctl_5_8)
        , .Y(\off_time[1] ));
    NOR3C \counter_RNIKM2J6[26]  (.A(\counter[25]_net_1 ), .B(
        counter_c24), .C(\counter[26]_net_1 ), .Y(counter_c26));
    NOR2A un1_counter_2_0_I_118 (.A(I_14_4), .B(\counter[5]_net_1 ), 
        .Y(N_14));
    OR2A un1_counter_0_I_103 (.A(\counter[14]_net_1 ), .B(
        \off_time[14] ), .Y(N_29));
    NOR2A \counter_RNO[28]  (.A(counter_n28_tz), .B(
        cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n28));
    XA1B \counter_RNO[15]  (.A(\counter[15]_net_1 ), .B(counter_c14), 
        .C(N_400_0), .Y(counter_n15));
    XNOR2 un1_counter_0_I_25 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .Y(\DWACT_BL_EQUAL_0_E_3[3] ));
    AND2 un1_counter_0_I_114 (.A(\DWACT_BL_EQUAL_0_E[4] ), .B(
        \DWACT_BL_EQUAL_0_E_0[3] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] ));
    XNOR2 un1_counter_0_I_11 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .Y(\DWACT_BL_EQUAL_0_E_4[3] ));
    OR3A un1_act_ctl_I_22 (.A(act_ctl_5_1), .B(\DWACT_FDEC_E[2] ), .C(
        \DWACT_FDEC_E[0] ), .Y(N_2_1));
    AX1C \counter_RNO_0[22]  (.A(\counter[21]_net_1 ), .B(counter_c20), 
        .C(\counter[22]_net_1 ), .Y(counter_n22_tz));
    XA1B \counter_RNO[7]  (.A(\counter[7]_net_1 ), .B(counter_c6), .C(
        N_400_0), .Y(counter_n7));
    OA1A un1_counter_2_0_I_125 (.A(N_16), .B(N_18), .C(N_17), .Y(N_21));
    DFN1E1C0 \off_reg[2]  (.D(off_div[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[2]_net_1 ));
    XNOR2 un1_counter_0_I_72 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .Y(\DWACT_BL_EQUAL_0_E_2[3] ));
    OA1 un1_counter_0_I_126 (.A(N_21_0), .B(N_20_0), .C(N_19), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] ));
    MX2C cur_pwm_RNIVKRSJ2_0 (.A(I_140_4), .B(I_140_3), .S(
        primary_fb_c), .Y(cur_pwm_RNIVKRSJ2_0_net_1));
    DFN1C0 \counter[6]  (.D(counter_n6), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[6]_net_1 ));
    AO1C un1_counter_0_I_122 (.A(\counter[7]_net_1 ), .B(\off_time[7] )
        , .C(N_12), .Y(N_18_0));
    XA1B \counter_RNO[31]  (.A(\counter[31]_net_1 ), .B(counter_63_0), 
        .C(cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n31));
    DFN1C0 \counter[21]  (.D(counter_n21), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[21]_net_1 ));
    AND2 un1_counter_0_I_20 (.A(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] ), .B(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] ), .Y(
        \DWACT_COMP0_E_0[1] ));
    OR2 un1_act_ctl_I_10 (.A(act_ctl_5), .B(act_ctl_5), .Y(
        \DWACT_FDEC_E[0] ));
    DFN1C0 \counter[3]  (.D(counter_n3), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[3]_net_1 ));
    DFN1C0 \counter[2]  (.D(counter_n2), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[2]_net_1 ));
    AND3 un1_counter_0_I_45 (.A(\DWACT_BL_EQUAL_0_E_3[2] ), .B(
        \DWACT_BL_EQUAL_0_E_2[1] ), .C(\DWACT_BL_EQUAL_0_E_3[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] ));
    DFN1E1C0 \off_reg[23]  (.D(off_div[23]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[23]_net_1 ));
    NOR2A \counter_RNO[8]  (.A(counter_n8_tz), .B(
        cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n8));
    OA1A un1_counter_2_0_I_121 (.A(\counter[8]_net_1 ), .B(I_23_6), .C(
        N_13), .Y(N_17));
    XA1B \counter_RNO[13]  (.A(\counter[13]_net_1 ), .B(counter_c12), 
        .C(N_400_0), .Y(counter_n13));
    NOR2B \counter_RNINUMD[13]  (.A(\counter[13]_net_1 ), .B(
        \counter[14]_net_1 ), .Y(counter_m6_0_a2_2));
    AO1C un1_counter_0_I_57 (.A(\off_time[20] ), .B(
        \counter[20]_net_1 ), .C(N_34), .Y(N_36));
    NOR3C \counter_RNI6PU12[5]  (.A(\counter[5]_net_1 ), .B(counter_c4)
        , .C(\counter[6]_net_1 ), .Y(counter_c6));
    DFN1E1C0 \off_reg[9]  (.D(off_div[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[9]_net_1 ));
    XNOR2 un1_counter_0_I_26 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(\DWACT_BL_EQUAL_0_E_4[2] ));
    AX1C \counter_RNO_0[4]  (.A(\counter[3]_net_1 ), .B(counter_c2), 
        .C(\counter[4]_net_1 ), .Y(counter_n4_tz));
    AO1C un1_counter_0_I_35 (.A(\off_time[28] ), .B(
        \counter[28]_net_1 ), .C(N_44), .Y(N_46));
    AO1 un1_counter_0_I_65 (.A(\DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] ), 
        .B(\DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] ), .C(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] ), .Y(\DWACT_COMP0_E[0] ));
    AND2 un1_counter_0_I_84 (.A(\DWACT_BL_EQUAL_0_E_1[3] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[1] ));
    NOR3C \counter_RNISENT1[11]  (.A(counter_m6_0_a2_2), .B(
        counter_m6_0_a2_1), .C(counter_m6_0_a2_6), .Y(
        counter_m6_0_a2_7));
    DFN1C0 cur_pwm (.D(cur_pwm_RNO_1), .CLK(clk_c), .CLR(n_rst_c), .Q(
        primary_fb_c));
    XA1B \counter_RNO[12]  (.A(\counter[12]_net_1 ), .B(counter_c11), 
        .C(N_400_0), .Y(counter_n12));
    NOR2A \off_reg_RNINT79[24]  (.A(\off_reg[24]_net_1 ), .B(
        act_ctl_5_2), .Y(\off_time[24] ));
    AOI1A un1_counter_0_I_95 (.A(\ACT_LT4_E[3] ), .B(\ACT_LT4_E[6] ), 
        .C(\ACT_LT4_E[10] ), .Y(\DWACT_CMPLE_PO0_DWACT_COMP0_E[0] ));
    OA1A un1_counter_0_I_40 (.A(N_46), .B(N_48), .C(N_47), .Y(N_51));
    XA1B \counter_RNO[1]  (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(N_400_0), .Y(counter_n1));
    DFN1C0 \counter[17]  (.D(counter_n17), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[17]_net_1 ));
    NOR2A \off_reg_RNIR189[28]  (.A(\off_reg[28]_net_1 ), .B(
        act_ctl_5_2), .Y(\off_time[28] ));
    NOR2 un1_counter_2_0_I_129 (.A(\counter[0]_net_1 ), .B(act_ctl_5_3)
        , .Y(N_4));
    DFN1C0 \counter[4]  (.D(counter_n4), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[4]_net_1 ));
    AO1B un1_counter_2_0_I_131 (.A(act_ctl_5_0), .B(\counter[1]_net_1 )
        , .C(N_4), .Y(N_6));
    NOR2B \counter_RNIG48E4[16]  (.A(counter_c15), .B(
        \counter[16]_net_1 ), .Y(counter_c16));
    AND2 un1_counter_0_I_30 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] ));
    OR2A un1_counter_0_I_60 (.A(\counter[23]_net_1 ), .B(
        \off_time[23] ), .Y(N_39));
    DFN1E1C0 \off_reg[11]  (.D(off_div[11]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[11]_net_1 ));
    AND2 un1_counter_0_I_29 (.A(\DWACT_BL_EQUAL_0_E_1[4] ), .B(
        \DWACT_BL_EQUAL_0_E_3[3] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] ));
    DFN1E1C0 \off_reg[22]  (.D(off_div[22]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[22]_net_1 ));
    DFN1C0 \counter[10]  (.D(counter_n10), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[10]_net_1 ));
    NOR2A un1_counter_2_0_I_19 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] ), .B(\counter[31]_net_1 )
        , .Y(\DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] ));
    NOR2A un1_counter_0_I_46 (.A(\off_time[24] ), .B(
        \counter[24]_net_1 ), .Y(\ACT_LT3_E[0] ));
    GND GND_i (.Y(GND));
    DFN1C0 \counter[13]  (.D(counter_n13), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[13]_net_1 ));
    XNOR2 un1_counter_0_I_81 (.A(\counter[16]_net_1 ), .B(
        \off_time[16] ), .Y(\DWACT_BL_EQUAL_0_E_0[1] ));
    NOR2A un1_counter_0_I_90 (.A(\off_time[18] ), .B(
        \counter[18]_net_1 ), .Y(\ACT_LT4_E[5] ));
    XNOR2 un1_counter_0_I_74 (.A(\counter[11]_net_1 ), .B(
        \off_time[11] ), .Y(\DWACT_BL_EQUAL_0_E_1[1] ));
    NOR2B un1_counter_2_0_I_140 (.A(\DWACT_COMP0_E[2] ), .B(
        \DWACT_COMP0_E[1] ), .Y(I_140_3));
    OA1A un1_counter_0_I_36 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .C(N_43), .Y(N_47));
    XNOR2 un1_counter_0_I_66 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\DWACT_BL_EQUAL_0_E[8] ));
    AND3 un1_counter_0_I_17 (.A(\DWACT_BL_EQUAL_0_E_5[0] ), .B(
        \DWACT_BL_EQUAL_0_E_4[1] ), .C(\DWACT_BL_EQUAL_0_E_5[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] ));
    DFN1E1C0 \off_reg[17]  (.D(off_div[17]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[17]_net_1 ));
    AX1C \counter_RNO_0[10]  (.A(\counter[9]_net_1 ), .B(counter_c8), 
        .C(\counter[10]_net_1 ), .Y(counter_n10_tz));
    DFN1C0 \counter[12]  (.D(counter_n12), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[12]_net_1 ));
    OR2A un1_counter_0_I_130 (.A(\off_time[4] ), .B(\counter[4]_net_1 )
        , .Y(N_5));
    NOR2B un1_counter_2_0_I_139 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E[2] )
        , .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ), .Y(
        \DWACT_COMP0_E[2] ));
    DFN1C0 \counter[27]  (.D(counter_n27), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[27]_net_1 ));
    OR2A un1_counter_0_I_96 (.A(\off_time[11] ), .B(
        \counter[11]_net_1 ), .Y(N_22));
    AOI1A un1_counter_0_I_49 (.A(\ACT_LT3_E[0] ), .B(\ACT_LT3_E[1] ), 
        .C(\ACT_LT3_E[2] ), .Y(\ACT_LT3_E[3] ));
    OR2 \off_reg_RNIR079[19]  (.A(\off_reg[19]_net_1 ), .B(act_ctl_5_2)
        , .Y(\off_time[19] ));
    AX1C \counter_RNO_0[20]  (.A(\counter[19]_net_1 ), .B(counter_c18), 
        .C(\counter[20]_net_1 ), .Y(counter_n20_tz));
    DFN1C0 \counter[20]  (.D(counter_n20), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[20]_net_1 ));
    OA1A un1_counter_0_I_101 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .C(N_23), .Y(N_27));
    DFN1E1C0 \off_reg[19]  (.D(off_div[19]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[19]_net_1 ));
    XNOR2 un1_counter_0_I_71 (.A(\counter[10]_net_1 ), .B(
        \off_time[10] ), .Y(\DWACT_BL_EQUAL_0_E_2[0] ));
    OR2A un1_counter_0_I_116 (.A(\off_time[6] ), .B(\counter[6]_net_1 )
        , .Y(N_12));
    AO1C un1_counter_0_I_39 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .C(N_45), .Y(N_50));
    XA1B \counter_RNO[17]  (.A(\counter[17]_net_1 ), .B(counter_c16), 
        .C(N_400_0), .Y(counter_n17));
    XNOR2 un1_counter_0_I_69 (.A(\counter[16]_net_1 ), .B(
        \off_time[16] ), .Y(\DWACT_BL_EQUAL_0_E[6] ));
    XNOR2 un1_counter_0_I_112 (.A(\counter[9]_net_1 ), .B(
        \off_time[9] ), .Y(\DWACT_BL_EQUAL_0_E[4] ));
    OA1A un1_counter_0_I_105 (.A(N_26), .B(N_28), .C(N_27), .Y(N_31));
    DFN1C0 \counter[23]  (.D(counter_n23), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[23]_net_1 ));
    NOR2A \off_reg_RNILR79[22]  (.A(\off_reg[22]_net_1 ), .B(
        act_ctl_5_2), .Y(\off_time[22] ));
    NOR3C \counter_RNIL1S07[27]  (.A(\counter[27]_net_1 ), .B(
        counter_c26), .C(\counter[28]_net_1 ), .Y(counter_c28));
    XA1B \counter_RNO[29]  (.A(\counter[29]_net_1 ), .B(counter_c28), 
        .C(cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n29));
    DFN1E1C0 \off_reg[25]  (.D(off_div[25]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[25]_net_1 ));
    NOR2B \counter_RNO_0[18]  (.A(counter_c16), .B(\counter[17]_net_1 )
        , .Y(counter_c17));
    DFN1C0 \counter[22]  (.D(counter_n22), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[22]_net_1 ));
    DFN1C0 \counter[15]  (.D(counter_n15), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[15]_net_1 ));
    AO1 un1_counter_0_I_107 (.A(\DWACT_CMPLE_PO0_DWACT_COMP0_E[1] ), 
        .B(\DWACT_CMPLE_PO0_DWACT_COMP0_E[2] ), .C(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] ));
    OR2A un1_counter_0_I_99 (.A(\off_time[14] ), .B(
        \counter[14]_net_1 ), .Y(N_25));
    NOR2A un1_counter_2_0_I_122 (.A(I_20_4), .B(\counter[7]_net_1 ), 
        .Y(N_18));
    AND2 un1_counter_2_0_I_115 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] ));
    XNOR2 un1_counter_0_I_108 (.A(\counter[5]_net_1 ), .B(
        \off_time[5] ), .Y(\DWACT_BL_EQUAL_0_E_0[0] ));
    NOR3C \counter_RNIFBVR4[9]  (.A(\counter[9]_net_1 ), .B(counter_c8)
        , .C(counter_m6_0_a2_7), .Y(counter_c18));
    AX1C \counter_RNO_0[8]  (.A(\counter[7]_net_1 ), .B(counter_c6), 
        .C(\counter[8]_net_1 ), .Y(counter_n8_tz));
    AX1C \counter_RNO_0[28]  (.A(\counter[27]_net_1 ), .B(counter_c26), 
        .C(\counter[28]_net_1 ), .Y(counter_n28_tz));
    VCC VCC_i (.Y(VCC));
    AO1C un1_counter_0_I_120 (.A(\off_time[6] ), .B(\counter[6]_net_1 )
        , .C(N_14_0), .Y(N_16_0));
    DFN1E1C0 \off_reg[31]  (.D(off_div[31]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[31]_net_1 ));
    XA1B \counter_RNO[14]  (.A(\counter[14]_net_1 ), .B(counter_c13), 
        .C(N_400_0), .Y(counter_n14));
    XNOR2 un1_counter_2_0_I_111 (.A(\counter[7]_net_1 ), .B(I_20_4), 
        .Y(\DWACT_BL_EQUAL_0_E[2] ));
    DFN1E1C0 \off_reg[7]  (.D(off_div[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[7]_net_1 ));
    DFN1C0 \counter[1]  (.D(counter_n1), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[1]_net_1 ));
    XNOR2 un1_counter_0_I_2 (.A(\counter[19]_net_1 ), .B(
        \off_time[19] ), .Y(\DWACT_BL_EQUAL_0_E_5[0] ));
    NOR2A \off_reg_RNIJP79[20]  (.A(\off_reg[20]_net_1 ), .B(
        act_ctl_5_2), .Y(\off_time[20] ));
    NOR2A \counter_RNO[26]  (.A(counter_n26_tz), .B(
        cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n26));
    NOR2A un1_counter_0_I_55 (.A(\off_time[19] ), .B(
        \counter[19]_net_1 ), .Y(N_34));
    AO1 un1_counter_0_I_139 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] ), .Y(\DWACT_COMP0_E_0[2] )
        );
    XA1B \counter_RNO[5]  (.A(\counter[5]_net_1 ), .B(counter_c4), .C(
        N_400_0), .Y(counter_n5));
    AO1C un1_counter_0_I_133 (.A(\counter[2]_net_1 ), .B(\off_time[2] )
        , .C(N_2_0), .Y(N_8_0));
    NOR2A \off_reg_RNICRPM[4]  (.A(\off_reg[4]_net_1 ), .B(act_ctl_5_9)
        , .Y(\off_time[4] ));
    DFN1C0 \counter[25]  (.D(counter_n25), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[25]_net_1 ));
    NOR2A \off_reg_RNIJM38[12]  (.A(\off_reg[12]_net_1 ), .B(
        act_ctl_5_1), .Y(\off_time[12] ));
    AND2A un1_counter_0_I_87 (.A(\off_time[16] ), .B(
        \counter[16]_net_1 ), .Y(\ACT_LT4_E[2] ));
    XA1B \counter_RNO[3]  (.A(\counter[3]_net_1 ), .B(counter_c2), .C(
        N_400_0), .Y(counter_n3));
    NOR2A \off_reg_RNIKQ79[21]  (.A(\off_reg[21]_net_1 ), .B(
        act_ctl_5_2), .Y(\off_time[21] ));
    DFN1E1C0 \off_reg[6]  (.D(off_div[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[6]_net_1 ));
    AND3 un1_counter_0_I_28 (.A(\DWACT_BL_EQUAL_0_E_4[0] ), .B(
        \DWACT_BL_EQUAL_0_E_3[1] ), .C(\DWACT_BL_EQUAL_0_E_4[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] ));
    NOR2A \off_reg_RNIMS79[23]  (.A(\off_reg[23]_net_1 ), .B(
        act_ctl_5_2), .Y(\off_time[23] ));
    OR2A un1_counter_0_I_50 (.A(\off_time[26] ), .B(
        \counter[26]_net_1 ), .Y(\ACT_LT3_E[4] ));
    DFN1C0 \counter[5]  (.D(counter_n5), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[5]_net_1 ));
    MX2A cur_pwm_RNO (.A(I_140_4), .B(I_140_3), .S(primary_fb_c), .Y(
        cur_pwm_RNO_1));
    XNOR2 un1_counter_0_I_4 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(\DWACT_BL_EQUAL_0_E[10] ));
    XNOR2 un1_counter_0_I_23 (.A(\counter[27]_net_1 ), .B(
        \off_time[27] ), .Y(\DWACT_BL_EQUAL_0_E_4[0] ));
    NOR2A \off_reg_RNILS89[31]  (.A(\off_reg[31]_net_1 ), .B(
        act_ctl_5_2), .Y(\off_time[31] ));
    NOR3C \counter_RNIIL921[18]  (.A(\counter[16]_net_1 ), .B(
        \counter[18]_net_1 ), .C(counter_m6_0_a2_4), .Y(
        counter_m6_0_a2_6));
    NOR2A \counter_RNO[10]  (.A(counter_n10_tz), .B(
        cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n10));
    AND3 un1_counter_0_I_77 (.A(\DWACT_BL_EQUAL_0_E_2[0] ), .B(
        \DWACT_BL_EQUAL_0_E_1[1] ), .C(\DWACT_BL_EQUAL_0_E_2[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] ));
    XNOR2 un1_counter_0_I_3 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .Y(\DWACT_BL_EQUAL_0_E[11] ));
    XA1B \counter_RNO[21]  (.A(\counter[21]_net_1 ), .B(counter_c20), 
        .C(N_400_0), .Y(counter_n21));
    XNOR2 un1_counter_0_I_6 (.A(\counter[20]_net_1 ), .B(
        \off_time[20] ), .Y(\DWACT_BL_EQUAL_0_E_4[1] ));
    OR2A un1_counter_0_I_56 (.A(\off_time[23] ), .B(
        \counter[23]_net_1 ), .Y(N_35));
    AX1C \counter_RNO_0[24]  (.A(\counter[23]_net_1 ), .B(counter_c22), 
        .C(\counter[24]_net_1 ), .Y(counter_n24_tz));
    AND3 un1_counter_0_I_15 (.A(\DWACT_BL_EQUAL_0_E_0[6] ), .B(
        \DWACT_BL_EQUAL_0_E_0[7] ), .C(\DWACT_BL_EQUAL_0_E_0[8] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] ));
    OR2 \off_reg_RNINQ38[16]  (.A(\off_reg[16]_net_1 ), .B(act_ctl_5_1)
        , .Y(\off_time[16] ));
    AND2A un1_counter_0_I_48 (.A(\off_time[25] ), .B(
        \counter[25]_net_1 ), .Y(\ACT_LT3_E[2] ));
    NOR2A un1_counter_0_I_129 (.A(\off_time[0] ), .B(
        \counter[0]_net_1 ), .Y(N_4_0));
    XNOR2 un1_counter_0_I_9 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(\DWACT_BL_EQUAL_0_E[12] ));
    AO1 un1_counter_0_I_140 (.A(\DWACT_COMP0_E_0[1] ), .B(
        \DWACT_COMP0_E_0[2] ), .C(\DWACT_COMP0_E[0] ), .Y(I_140_4));
    OR2A un1_counter_0_I_123 (.A(\counter[9]_net_1 ), .B(\off_time[9] )
        , .Y(N_19));
    DFN1C0 \counter[16]  (.D(counter_n16), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[16]_net_1 ));
    OR2A un1_counter_0_I_38 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(N_49));
    OR2 \off_reg_RNIH0QM[9]  (.A(\off_reg[9]_net_1 ), .B(act_ctl_5_9), 
        .Y(\off_time[9] ));
    XA1B \counter_RNO[25]  (.A(\counter[25]_net_1 ), .B(counter_c24), 
        .C(cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n25));
    XNOR2 un1_counter_0_I_68 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\DWACT_BL_EQUAL_0_E[7] ));
    NOR3C \counter_RNIOD8S[2]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .C(\counter[2]_net_1 ), .Y(counter_c2));
    XNOR2 un1_act_ctl_I_14 (.A(N_5_0), .B(act_ctl_5), .Y(I_14_4));
    NOR2B \counter_RNO_0[31]  (.A(\counter[30]_net_1 ), .B(counter_c29)
        , .Y(counter_63_0));
    XNOR2 un1_counter_0_I_43 (.A(\counter[25]_net_1 ), .B(
        \off_time[25] ), .Y(\DWACT_BL_EQUAL_0_E_2[1] ));
    XOR2 un1_act_ctl_I_20 (.A(act_ctl_5), .B(N_3), .Y(I_20_4));
    AO1C un1_counter_0_I_59 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .C(N_32), .Y(N_38));
    DFN1E1C0 \off_reg[21]  (.D(off_div[21]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[21]_net_1 ));
    AO1C un1_counter_0_I_104 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .C(N_25), .Y(N_30));
    OR2 un1_counter_2_0_I_127 (.A(\counter[1]_net_1 ), .B(act_ctl_5_3), 
        .Y(N_2));
    XNOR2 un1_counter_0_I_10 (.A(\counter[24]_net_1 ), .B(
        \off_time[24] ), .Y(\DWACT_BL_EQUAL_0_E_0[5] ));
    NOR2A un1_counter_0_I_98 (.A(\off_time[10] ), .B(
        \counter[10]_net_1 ), .Y(N_24));
    NOR2A un1_counter_0_I_33 (.A(\off_time[27] ), .B(
        \counter[27]_net_1 ), .Y(N_44));
    OA1 un1_counter_0_I_63 (.A(N_41), .B(N_40), .C(N_39), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] ));
    NOR2A \counter_RNO[6]  (.A(counter_n6_tz), .B(
        cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n6));
    XA1B \counter_RNO[30]  (.A(\counter[30]_net_1 ), .B(counter_c29), 
        .C(cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n30));
    NOR2A \off_reg_RNIOU79[25]  (.A(\off_reg[25]_net_1 ), .B(
        act_ctl_5_2), .Y(\off_time[25] ));
    OR2 \off_reg_RNIQV69[18]  (.A(\off_reg[18]_net_1 ), .B(act_ctl_5_2)
        , .Y(\off_time[18] ));
    XNOR2 un1_counter_0_I_110 (.A(\counter[8]_net_1 ), .B(
        \off_time[8] ), .Y(\DWACT_BL_EQUAL_0_E_0[3] ));
    DFN1E1C0 \off_reg[27]  (.D(off_div[27]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[27]_net_1 ));
    AND3 un1_counter_0_I_16 (.A(\DWACT_BL_EQUAL_0_E_4[3] ), .B(
        \DWACT_BL_EQUAL_0_E_2[4] ), .C(\DWACT_BL_EQUAL_0_E_0[5] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] ));
    OR2A un1_counter_0_I_93 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\ACT_LT4_E[8] ));
    DFN1E1C0 \off_reg[8]  (.D(off_div[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[8]_net_1 ));
    DFN1C0 \counter[26]  (.D(counter_n26), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[26]_net_1 ));
    XA1B \counter_RNO[23]  (.A(\counter[23]_net_1 ), .B(counter_c22), 
        .C(N_400_0), .Y(counter_n23));
    NOR2A \off_reg_RNIKN38[13]  (.A(\off_reg[13]_net_1 ), .B(
        act_ctl_5_1), .Y(\off_time[13] ));
    NOR2A \off_reg_RNI7KML[0]  (.A(\off_reg[0]_net_1 ), .B(act_ctl_5_8)
        , .Y(\off_time[0] ));
    OA1C un1_counter_2_0_I_137 (.A(\counter[3]_net_1 ), .B(N_11), .C(
        \counter[4]_net_1 ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] ));
    OR2B un1_counter_2_0_I_133 (.A(N_2), .B(\counter[2]_net_1 ), .Y(
        N_8));
    OR2 un1_act_ctl_I_19 (.A(\DWACT_FDEC_E[2] ), .B(\DWACT_FDEC_E[0] ), 
        .Y(N_3));
    DFN1C0 \counter[14]  (.D(counter_n14), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[14]_net_1 ));
    DFN1E1C0 \off_reg[29]  (.D(off_div[29]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[29]_net_1 ));
    AND3 un1_counter_2_0_I_18 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] ));
    DFN1E1C0 \off_reg[1]  (.D(off_div[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[1]_net_1 ));
    NOR2A \counter_RNO[22]  (.A(counter_n22_tz), .B(
        cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n22));
    AO1C un1_counter_0_I_131 (.A(\off_time[1] ), .B(\counter[1]_net_1 )
        , .C(N_4_0), .Y(N_6_0));
    AND2 un1_counter_0_I_19 (.A(\DWACT_BL_EQUAL_0_E[12] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] ));
    XNOR2 un1_counter_0_I_42 (.A(\counter[26]_net_1 ), .B(
        \off_time[26] ), .Y(\DWACT_BL_EQUAL_0_E_3[2] ));
    AO1C un1_counter_0_I_135 (.A(\counter[3]_net_1 ), .B(\off_time[3] )
        , .C(N_5), .Y(N_10));
    DFN1E1C0 \off_reg[10]  (.D(off_div[10]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[10]_net_1 ));
    NOR2A un1_counter_0_I_85 (.A(\off_time[15] ), .B(
        \counter[15]_net_1 ), .Y(\ACT_LT4_E[0] ));
    DFN1C0 \counter[31]  (.D(counter_n31), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[31]_net_1 ));
    OR2A un1_counter_0_I_32 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(N_43));
    OA1A un1_counter_0_I_62 (.A(N_36), .B(N_38), .C(N_37), .Y(N_41));
    OR3A un1_act_ctl_I_13 (.A(act_ctl_5_1), .B(act_ctl_5_1), .C(
        \DWACT_FDEC_E[0] ), .Y(N_5_0));
    OA1 un1_counter_0_I_137 (.A(N_11_0), .B(N_10), .C(N_9), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] ));
    NOR3C \counter_RNIUCGN5[22]  (.A(\counter[21]_net_1 ), .B(
        counter_c20), .C(\counter[22]_net_1 ), .Y(counter_c22));
    NOR3C \counter_RNIDH3F1[4]  (.A(\counter[3]_net_1 ), .B(counter_c2)
        , .C(\counter[4]_net_1 ), .Y(counter_c4));
    AO1 un1_counter_0_I_138 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] ));
    NOR2A un1_counter_0_I_92 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\ACT_LT4_E[7] ));
    DFN1C0 \counter[24]  (.D(counter_n24), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[24]_net_1 ));
    OR2A un1_counter_0_I_119 (.A(\off_time[9] ), .B(\counter[9]_net_1 )
        , .Y(N_15));
    NOR3 un1_counter_2_0_I_14 (.A(\counter[29]_net_1 ), .B(
        \counter[30]_net_1 ), .C(\counter[28]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] ));
    AND3 un1_counter_2_0_I_78 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ));
    XNOR2 un1_counter_0_I_80 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\DWACT_BL_EQUAL_0_E_1[2] ));
    XNOR2 un1_counter_0_I_5 (.A(\counter[27]_net_1 ), .B(
        \off_time[27] ), .Y(\DWACT_BL_EQUAL_0_E_0[8] ));
    AND3 un1_counter_0_I_113 (.A(\DWACT_BL_EQUAL_0_E_0[0] ), .B(
        \DWACT_BL_EQUAL_0_E[1] ), .C(\DWACT_BL_EQUAL_0_E_0[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] ));
    XNOR2 un1_counter_0_I_24 (.A(\counter[28]_net_1 ), .B(
        \off_time[28] ), .Y(\DWACT_BL_EQUAL_0_E_3[1] ));
    NOR2A \counter_RNO[4]  (.A(counter_n4_tz), .B(
        cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n4));
    AND3 un1_counter_0_I_75 (.A(\DWACT_BL_EQUAL_0_E[6] ), .B(
        \DWACT_BL_EQUAL_0_E[7] ), .C(\DWACT_BL_EQUAL_0_E[8] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] ));
    DFN1E1C0 \off_reg[14]  (.D(off_div[14]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[14]_net_1 ));
    NOR3C \counter_RNI35QK2[8]  (.A(\counter[7]_net_1 ), .B(counter_c6)
        , .C(\counter[8]_net_1 ), .Y(counter_c8));
    NOR2A \off_reg_RNIPV79[26]  (.A(\off_reg[26]_net_1 ), .B(
        act_ctl_5_2), .Y(\off_time[26] ));
    NOR2A \off_reg_RNIFUPM[7]  (.A(\off_reg[7]_net_1 ), .B(act_ctl_5_9)
        , .Y(\off_time[7] ));
    OR2A un1_counter_2_0_I_120 (.A(N_14), .B(\counter[6]_net_1 ), .Y(
        N_16));
    XA1B \counter_RNO[18]  (.A(\counter[18]_net_1 ), .B(counter_c17), 
        .C(N_400_0), .Y(counter_n18));
    NOR3 un1_counter_2_0_I_15 (.A(\counter[26]_net_1 ), .B(
        \counter[27]_net_1 ), .C(\counter[25]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] ));
    OR2A un1_counter_0_I_86 (.A(\off_time[16] ), .B(
        \counter[16]_net_1 ), .Y(\ACT_LT4_E[1] ));
    NOR2A un1_counter_2_0_I_124 (.A(I_23_6), .B(\counter[8]_net_1 ), 
        .Y(N_20));
    OA1A un1_counter_0_I_58 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .C(N_33), .Y(N_37));
    OA1A un1_counter_0_I_121 (.A(\counter[8]_net_1 ), .B(\off_time[8] )
        , .C(N_13_0), .Y(N_17_0));
    AND2 un1_counter_2_0_I_20 (.A(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] ), .B(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] ), .Y(
        \DWACT_COMP0_E[1] ));
    AX1C \counter_RNO_0[26]  (.A(\counter[25]_net_1 ), .B(counter_c24), 
        .C(\counter[26]_net_1 ), .Y(counter_n26_tz));
    XA1B \counter_RNO[27]  (.A(\counter[27]_net_1 ), .B(counter_c26), 
        .C(cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n27));
    NOR2A \off_reg_RNIGVPM[8]  (.A(\off_reg[8]_net_1 ), .B(act_ctl_5_9)
        , .Y(\off_time[8] ));
    OA1A un1_counter_0_I_125 (.A(N_16_0), .B(N_18_0), .C(N_17_0), .Y(
        N_21_0));
    AX1C \counter_RNO_0[6]  (.A(\counter[5]_net_1 ), .B(counter_c4), 
        .C(\counter[6]_net_1 ), .Y(counter_n6_tz));
    XNOR2 un1_counter_0_I_70 (.A(\counter[15]_net_1 ), .B(
        \off_time[15] ), .Y(\DWACT_BL_EQUAL_0_E[5] ));
    OA1 un1_counter_0_I_106 (.A(N_31), .B(N_30), .C(N_29), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] ));
    DFN1E1C0 \off_reg[18]  (.D(off_div[18]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[18]_net_1 ));
    NOR2B \counter_RNIU2QI3[12]  (.A(counter_c11), .B(
        \counter[12]_net_1 ), .Y(counter_c12));
    AO1C un1_counter_0_I_102 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .C(N_22), .Y(N_28));
    OR2A un1_counter_2_0_I_117 (.A(\counter[7]_net_1 ), .B(I_20_4), .Y(
        N_13));
    NOR3B un1_counter_2_0_I_113 (.A(\DWACT_BL_EQUAL_0_E[2] ), .B(
        \DWACT_BL_EQUAL_0_E[0] ), .C(\counter[6]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ));
    XNOR2 un1_counter_0_I_44 (.A(\counter[24]_net_1 ), .B(
        \off_time[24] ), .Y(\DWACT_BL_EQUAL_0_E_3[0] ));
    OR2A un1_counter_0_I_53 (.A(\off_time[20] ), .B(
        \counter[20]_net_1 ), .Y(N_32));
    OR2A un1_counter_0_I_127 (.A(\off_time[1] ), .B(\counter[1]_net_1 )
        , .Y(N_2_0));
    MX2C cur_pwm_RNIVKRSJ2 (.A(I_140_4), .B(I_140_3), .S(primary_fb_c), 
        .Y(N_400_0));
    NOR2B \counter_RNIIIC74[15]  (.A(counter_c14), .B(
        \counter[15]_net_1 ), .Y(counter_c15));
    OR2A un1_counter_0_I_34 (.A(\off_time[31] ), .B(
        \counter[31]_net_1 ), .Y(N_45));
    OR2A un1_counter_0_I_128 (.A(\counter[2]_net_1 ), .B(\off_time[2] )
        , .Y(N_3_0));
    OR2A un1_counter_0_I_89 (.A(\off_time[17] ), .B(
        \counter[17]_net_1 ), .Y(\ACT_LT4_E[4] ));
    AO1 un1_counter_0_I_64 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] ));
    DFN1E1C0 \off_reg[16]  (.D(off_div[16]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[16]_net_1 ));
    AND3 un1_counter_0_I_76 (.A(\DWACT_BL_EQUAL_0_E_2[3] ), .B(
        \DWACT_BL_EQUAL_0_E_0[4] ), .C(\DWACT_BL_EQUAL_0_E[5] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] ));
    XNOR2 un1_counter_0_I_1 (.A(\counter[23]_net_1 ), .B(
        \off_time[23] ), .Y(\DWACT_BL_EQUAL_0_E_2[4] ));
    DFN1E1C0 \off_reg[30]  (.D(off_div[30]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[30]_net_1 ));
    NOR3 un1_counter_2_0_I_75 (.A(\counter[17]_net_1 ), .B(
        \counter[18]_net_1 ), .C(\counter[16]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] ));
    NOR2A \counter_RNO[24]  (.A(counter_n24_tz), .B(
        cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n24));
    DFN1C0 \counter[7]  (.D(counter_n7), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[7]_net_1 ));
    AOI1A un1_counter_0_I_94 (.A(\ACT_LT4_E[7] ), .B(\ACT_LT4_E[8] ), 
        .C(\ACT_LT4_E[5] ), .Y(\ACT_LT4_E[10] ));
    DFN1C0 \counter[30]  (.D(counter_n30), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[30]_net_1 ));
    OA1 un1_counter_0_I_41 (.A(N_51), .B(N_50), .C(N_49), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] ));
    AND3 un1_counter_0_I_18 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] ));
    NOR2B \counter_RNINOO77[29]  (.A(counter_c28), .B(
        \counter[29]_net_1 ), .Y(counter_c29));
    OR2A un1_counter_0_I_31 (.A(\off_time[28] ), .B(
        \counter[28]_net_1 ), .Y(N_42));
    NOR2A \off_reg_RNIIL38[11]  (.A(\off_reg[11]_net_1 ), .B(
        act_ctl_5_1), .Y(\off_time[11] ));
    XNOR2 un1_counter_2_0_I_108 (.A(\counter[5]_net_1 ), .B(I_14_4), 
        .Y(\DWACT_BL_EQUAL_0_E[0] ));
    AO1C un1_counter_0_I_61 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .C(N_35), .Y(N_40));
    NOR2 \counter_RNO[0]  (.A(\counter[0]_net_1 ), .B(
        cur_pwm_RNIVKRSJ2_0_net_1), .Y(\counter_RNO_1[0] ));
    NOR3C \counter_RNIKFIK[10]  (.A(\counter[15]_net_1 ), .B(
        \counter[10]_net_1 ), .C(\counter[17]_net_1 ), .Y(
        counter_m6_0_a2_4));
    XNOR2 un1_counter_0_I_79 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\DWACT_BL_EQUAL_0_E_1[3] ));
    NOR2A \off_reg_RNIHK38[10]  (.A(\off_reg[10]_net_1 ), .B(
        act_ctl_5_1), .Y(\off_time[10] ));
    DFN1E1C0 \off_reg[3]  (.D(off_div[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[3]_net_1 ));
    NOR2B \counter_RNIJQMD[11]  (.A(\counter[11]_net_1 ), .B(
        \counter[12]_net_1 ), .Y(counter_m6_0_a2_1));
    DFN1E1C0 \off_reg[0]  (.D(off_div[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[0]_net_1 ));
    OR3 un1_act_ctl_I_18 (.A(act_ctl_5_1), .B(act_ctl_5_i), .C(
        act_ctl_5_1), .Y(\DWACT_FDEC_E[2] ));
    NOR2A \off_reg_RNIANML[3]  (.A(\off_reg[3]_net_1 ), .B(act_ctl_5_8)
        , .Y(\off_time[3] ));
    NOR2B \counter_RNIL1H04[14]  (.A(counter_c13), .B(
        \counter[14]_net_1 ), .Y(counter_c14));
    OA1B un1_counter_2_0_I_126 (.A(N_20), .B(N_21), .C(
        \counter[9]_net_1 ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ));
    OR2A un1_counter_0_I_134 (.A(\counter[4]_net_1 ), .B(\off_time[4] )
        , .Y(N_9));
    XNOR2 un1_counter_0_I_13 (.A(\counter[28]_net_1 ), .B(
        \off_time[28] ), .Y(\DWACT_BL_EQUAL_0_E[9] ));
    NOR2A un1_counter_0_I_91 (.A(\ACT_LT4_E[4] ), .B(\ACT_LT4_E[5] ), 
        .Y(\ACT_LT4_E[6] ));
    AOI1A un1_counter_0_I_52 (.A(\ACT_LT3_E[3] ), .B(\ACT_LT3_E[4] ), 
        .C(\ACT_LT3_E[5] ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] ));
    OR2 \off_reg_RNIETPM[6]  (.A(\off_reg[6]_net_1 ), .B(act_ctl_5_9), 
        .Y(\off_time[6] ));
    NOR2A \counter_RNO[20]  (.A(counter_n20_tz), .B(
        cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n20));
    DFN1E1C0 \off_reg[13]  (.D(off_div[13]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[13]_net_1 ));
    XNOR2 un1_counter_0_I_27 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(\DWACT_BL_EQUAL_0_E_1[4] ));
    XNOR2 un1_counter_0_I_111 (.A(\counter[7]_net_1 ), .B(
        \off_time[7] ), .Y(\DWACT_BL_EQUAL_0_E_0[2] ));
    OR2A un1_counter_2_0_I_136 (.A(N_6), .B(N_8), .Y(N_11));
    NOR2B \counter_RNI4LUB3[11]  (.A(counter_c10), .B(
        \counter[11]_net_1 ), .Y(counter_c11));
    OR2 \off_reg_RNIOR38[17]  (.A(\off_reg[17]_net_1 ), .B(act_ctl_5_1)
        , .Y(\off_time[17] ));
    AND2 un1_counter_0_I_115 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] ));
    DFN1E1C0 \off_reg[4]  (.D(off_div[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[4]_net_1 ));
    NOR3C \counter_RNIB8353[10]  (.A(\counter[9]_net_1 ), .B(
        counter_c8), .C(\counter[10]_net_1 ), .Y(counter_c10));
    XNOR2 un1_counter_2_0_I_110 (.A(\counter[8]_net_1 ), .B(I_23_6), 
        .Y(\DWACT_BL_EQUAL_0_E[3] ));
    XNOR2 un1_counter_0_I_8 (.A(\counter[25]_net_1 ), .B(
        \off_time[25] ), .Y(\DWACT_BL_EQUAL_0_E_0[6] ));
    DFN1E1C0 \off_reg[20]  (.D(off_div[20]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[20]_net_1 ));
    NOR2A \counter_RNO[2]  (.A(counter_n2_tz), .B(
        cur_pwm_RNIVKRSJ2_0_net_1), .Y(counter_n2));
    DFN1C0 \counter[9]  (.D(counter_n9), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[9]_net_1 ));
    NOR3 un1_counter_2_0_I_16 (.A(\counter[24]_net_1 ), .B(
        \counter[23]_net_1 ), .C(\counter[22]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] ));
    NOR2A un1_counter_2_0_I_114 (.A(\DWACT_BL_EQUAL_0_E[3] ), .B(
        \counter[9]_net_1 ), .Y(\DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ));
    OR2A un1_counter_0_I_117 (.A(\counter[7]_net_1 ), .B(\off_time[7] )
        , .Y(N_13_0));
    NOR3C \counter_RNINF956[24]  (.A(\counter[23]_net_1 ), .B(
        counter_c22), .C(\counter[24]_net_1 ), .Y(counter_c24));
    XA1B \counter_RNO[19]  (.A(\counter[19]_net_1 ), .B(counter_c18), 
        .C(N_400_0), .Y(counter_n19));
    AO1C un1_counter_0_I_124 (.A(\counter[8]_net_1 ), .B(\off_time[8] )
        , .C(N_15), .Y(N_20_0));
    NOR2A un1_counter_0_I_118 (.A(\off_time[5] ), .B(
        \counter[5]_net_1 ), .Y(N_14_0));
    XNOR2 un1_counter_0_I_12 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .Y(\DWACT_BL_EQUAL_0_E_5[2] ));
    AO1 un1_counter_2_0_I_138 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] )
        , .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] ));
    XA1B \counter_RNO[9]  (.A(\counter[9]_net_1 ), .B(counter_c8), .C(
        N_400_0), .Y(counter_n9));
    DFN1E1C0 \off_reg[12]  (.D(off_div[12]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[12]_net_1 ));
    AOI1A un1_counter_0_I_88 (.A(\ACT_LT4_E[0] ), .B(\ACT_LT4_E[1] ), 
        .C(\ACT_LT4_E[2] ), .Y(\ACT_LT4_E[3] ));
    OR2A un1_counter_0_I_47 (.A(\off_time[25] ), .B(
        \counter[25]_net_1 ), .Y(\ACT_LT3_E[1] ));
    NOR2A \off_reg_RNIKR89[30]  (.A(\off_reg[30]_net_1 ), .B(
        act_ctl_5_2), .Y(\off_time[30] ));
    DFN1C0 \counter[8]  (.D(counter_n8), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[8]_net_1 ));
    OR2A un1_counter_0_I_54 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .Y(N_33));
    AO1C un1_counter_0_I_37 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .C(N_42), .Y(N_48));
    XNOR2 un1_counter_0_I_7 (.A(\counter[26]_net_1 ), .B(
        \off_time[26] ), .Y(\DWACT_BL_EQUAL_0_E_0[7] ));
    XNOR2 un1_counter_0_I_67 (.A(\counter[14]_net_1 ), .B(
        \off_time[14] ), .Y(\DWACT_BL_EQUAL_0_E_0[4] ));
    DFN1C0 \counter[18]  (.D(counter_n18), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[18]_net_1 ));
    AO1C un1_counter_0_I_100 (.A(\off_time[11] ), .B(
        \counter[11]_net_1 ), .C(N_24), .Y(N_26));
    NOR2B \counter_RNIPHLP3[13]  (.A(counter_c12), .B(
        \counter[13]_net_1 ), .Y(counter_c13));
    DFN1E1C0 \off_reg[24]  (.D(off_div[24]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[24]_net_1 ));
    AND3 un1_counter_0_I_83 (.A(\DWACT_BL_EQUAL_0_E_1[0] ), .B(
        \DWACT_BL_EQUAL_0_E_0[1] ), .C(\DWACT_BL_EQUAL_0_E_1[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] ));
    XA1B \counter_RNO[16]  (.A(\counter[16]_net_1 ), .B(counter_c15), 
        .C(N_400_0), .Y(counter_n16));
    DFN1C0 \counter[0]  (.D(\counter_RNO_1[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\counter[0]_net_1 ));
    NOR3 un1_counter_2_0_I_76 (.A(\counter[15]_net_1 ), .B(
        \counter[14]_net_1 ), .C(\counter[13]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] ));
    OR2A un1_counter_0_I_97 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .Y(N_23));
    OR2 \off_reg_RNILO38[14]  (.A(\off_reg[14]_net_1 ), .B(act_ctl_5_1)
        , .Y(\off_time[14] ));
    
endmodule


module spi_clk_11s_3_0(
       sck_33_c,
       n_rst_c,
       clk_c
    );
output sck_33_c;
input  n_rst_c;
input  clk_c;

    wire N_8, \counter[1]_net_1 , \counter[0]_net_1 , N_6, 
        \counter[3]_net_1 , \DWACT_FINC_E[0] , cur_clk5_5, cur_clk5_3, 
        \counter[6]_net_1 , cur_clk5_4, cur_clk5_1, \counter[7]_net_1 , 
        \counter[8]_net_1 , \counter[4]_net_1 , \counter[5]_net_1 , 
        \counter[2]_net_1 , cur_clk_RNO_1, \counter_3[1] , I_5_1, 
        \counter_3[0] , \counter_3[3] , I_9_1, I_7_1, I_12_2, I_14_3, 
        I_17_2, I_20_3, I_23_4, N_2, \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[3] , N_3, N_4, \DWACT_FINC_E[1] , N_5, N_7, GND, 
        VCC;
    
    NOR2B un3_counter_I_6 (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(N_8));
    AND3 un3_counter_I_19 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\counter[6]_net_1 ), .Y(N_3));
    XOR2 un3_counter_I_20 (.A(N_3), .B(\counter[7]_net_1 ), .Y(I_20_3));
    DFN1C0 \counter[2]  (.D(I_7_1), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[2]_net_1 ));
    NOR2 \counter_RNI382P[2]  (.A(\counter[5]_net_1 ), .B(
        \counter[2]_net_1 ), .Y(cur_clk5_1));
    DFN1C0 \counter[7]  (.D(I_20_3), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[7]_net_1 ));
    AND3 un3_counter_I_13 (.A(\DWACT_FINC_E[0] ), .B(
        \counter[3]_net_1 ), .C(\counter[4]_net_1 ), .Y(N_5));
    AOI1 \counter_RNO[0]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(
        \counter[0]_net_1 ), .Y(\counter_3[0] ));
    DFN1C0 \counter[6]  (.D(I_17_2), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[6]_net_1 ));
    VCC VCC_i (.Y(VCC));
    XOR2 un3_counter_I_12 (.A(N_6), .B(\counter[4]_net_1 ), .Y(I_12_2));
    DFN1C0 \counter[8]  (.D(I_23_4), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[8]_net_1 ));
    NOR3A \counter_RNIEO4I1[8]  (.A(cur_clk5_1), .B(\counter[7]_net_1 )
        , .C(\counter[8]_net_1 ), .Y(cur_clk5_4));
    XOR2 un3_counter_I_23 (.A(N_2), .B(\counter[8]_net_1 ), .Y(I_23_4));
    AOI1B \counter_RNO[1]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(I_5_1), 
        .Y(\counter_3[1] ));
    AND3 un3_counter_I_22 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\DWACT_FINC_E[3] ), .Y(N_2));
    XOR2 un3_counter_I_7 (.A(N_8), .B(\counter[2]_net_1 ), .Y(I_7_1));
    NOR2B un3_counter_I_11 (.A(\counter[3]_net_1 ), .B(
        \DWACT_FINC_E[0] ), .Y(N_6));
    AND3 un3_counter_I_16 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[1] )
        , .C(\counter[5]_net_1 ), .Y(N_4));
    DFN1C0 \counter[4]  (.D(I_12_2), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[4]_net_1 ));
    XOR2 un3_counter_I_17 (.A(N_4), .B(\counter[6]_net_1 ), .Y(I_17_2));
    DFN1C0 \counter[5]  (.D(I_14_3), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[5]_net_1 ));
    AND3 un3_counter_I_8 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(N_7));
    GND GND_i (.Y(GND));
    AX1C cur_clk_RNO (.A(cur_clk5_4), .B(cur_clk5_5), .C(sck_33_c), .Y(
        cur_clk_RNO_1));
    AOI1B \counter_RNO[3]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(I_9_1), 
        .Y(\counter_3[3] ));
    AND2 un3_counter_I_21 (.A(\counter[6]_net_1 ), .B(
        \counter[7]_net_1 ), .Y(\DWACT_FINC_E[3] ));
    DFN1C0 \counter[1]  (.D(\counter_3[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[1]_net_1 ));
    NOR2A \counter_RNI382P[4]  (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(cur_clk5_3));
    DFN1C0 \counter[3]  (.D(\counter_3[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[3]_net_1 ));
    NOR3B \counter_RNI6G4I1[6]  (.A(\counter[1]_net_1 ), .B(cur_clk5_3)
        , .C(\counter[6]_net_1 ), .Y(cur_clk5_5));
    AND2 un3_counter_I_15 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(\DWACT_FINC_E[1] ));
    XOR2 un3_counter_I_9 (.A(N_7), .B(\counter[3]_net_1 ), .Y(I_9_1));
    DFN1C0 cur_clk (.D(cur_clk_RNO_1), .CLK(clk_c), .CLR(n_rst_c), .Q(
        sck_33_c));
    XOR2 un3_counter_I_14 (.A(N_5), .B(\counter[5]_net_1 ), .Y(I_14_3));
    XOR2 un3_counter_I_5 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .Y(I_5_1));
    AND3 un3_counter_I_10 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(
        \DWACT_FINC_E[0] ));
    DFN1C0 \counter[0]  (.D(\counter_3[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[0]_net_1 ));
    AND3 un3_counter_I_18 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .C(\counter[5]_net_1 ), .Y(
        \DWACT_FINC_E[2] ));
    
endmodule


module PID_controller_Z3_0(
       LED_12_0,
       LED_15_0,
       choose_0_0,
       LED_c_0,
       LED_5_0,
       choose,
       LED_33_0,
       LED_FB,
       primary_fb_c,
       act_ctl_5,
       act_ctl_5_8,
       act_ctl_5_9,
       act_ctl_5_1,
       act_ctl_5_2,
       act_ctl_5_0,
       act_ctl_5_3,
       act_ctl_5_i,
       din_fb_c,
       cs_i_1_i,
       sck_33_c,
       clk_c,
       n_rst_c
    );
input  LED_12_0;
input  LED_15_0;
input  choose_0_0;
output LED_c_0;
input  LED_5_0;
input  [2:0] choose;
input  LED_33_0;
output [7:0] LED_FB;
output primary_fb_c;
input  act_ctl_5;
input  act_ctl_5_8;
input  act_ctl_5_9;
input  act_ctl_5_1;
input  act_ctl_5_2;
input  act_ctl_5_0;
input  act_ctl_5_3;
input  act_ctl_5_i;
input  din_fb_c;
output cs_i_1_i;
output sck_33_c;
input  clk_c;
input  n_rst_c;

    wire \state[1] , \state[0] , pwm_chg, int_done, sig_prev, 
        sig_old_i_0, avg_done, int_enable, vd_rdy, sum_rdy, 
        deriv_enable, calc_avg, calc_int, pwm_enable, sum_enable, 
        avg_enable, pwm_chg_0, int_enable_0, int_enable_1, 
        int_enable_2, int_enable_3, int_enable_4, int_enable_5, 
        int_enable_6, int_enable_7, int_enable_8, int_enable_9, 
        int_enable_10, int_enable_11, int_enable_12, int_enable_13, 
        int_enable_14, int_enable_15, int_enable_16, int_enable_17, 
        int_enable_18, int_enable_19, int_enable_20, int_enable_21, 
        int_enable_22, int_enable_23, int_enable_24, int_enable_25, 
        int_enable_26, int_enable_27, int_enable_28, int_enable_29, 
        int_enable_30, int_enable_31, int_enable_32, int_enable_33, 
        avg_enable_0, avg_enable_1, calc_error, \cur_vd[0] , 
        \cur_vd[1] , \cur_vd[2] , \cur_vd[3] , \cur_vd[4] , 
        \cur_vd[5] , \cur_vd[6] , \cur_vd[7] , \cur_vd[8] , 
        \cur_vd[9] , \cur_vd[10] , \cur_vd[11] , \avg_new[0] , 
        \avg_new[1] , \avg_new[2] , \avg_new[3] , \avg_new[4] , 
        \avg_new[5] , \avg_new[6] , \avg_new[7] , \avg_new[8] , 
        \avg_new[9] , \avg_new[10] , \avg_new[11] , \avg_old[0] , 
        \avg_old[1] , \avg_old[2] , \avg_old[3] , \avg_old[4] , 
        \avg_old[5] , \avg_old[6] , \avg_old[7] , \avg_old[8] , 
        \avg_old[9] , \avg_old[10] , \avg_old[11] , \cur_error[0] , 
        \cur_error[1] , \cur_error[2] , \cur_error[3] , \cur_error[4] , 
        \cur_error[5] , \cur_error[6] , \cur_error[7] , \cur_error[8] , 
        \cur_error[9] , \cur_error[10] , \cur_error[11] , 
        \cur_error[12] , \LED_FB_i[5] , \LED_FB[4] , \average[2] , 
        \average[3] , \average[4] , \average[5] , \average[6] , 
        \sr_old[0] , \sr_old[1] , \sr_old[2] , \sr_old[3] , 
        \sr_old[4] , \sr_old[5] , \sr_old[6] , \sr_old[7] , 
        \sr_old[8] , \sr_old[9] , \sr_old[10] , \sr_old[11] , 
        \sr_old[12] , \sr_new[0] , \sr_new[1] , \sr_new[2] , 
        \sr_new[3] , \sr_new[4] , \sr_new[5] , \sr_new[6] , 
        \sr_new[7] , \sr_new[8] , \sr_new[9] , \sr_new[10] , 
        \sr_new[11] , \sr_new[12] , \sr_prev[0] , \sr_prev[1] , 
        \sr_prev[2] , \sr_prev[3] , \sr_prev[4] , \sr_prev[5] , 
        \sr_prev[6] , \sr_prev[7] , \sr_prev[8] , \sr_prev[9] , 
        \sr_prev[10] , \sr_prev[11] , \sr_prev[12] , \sr_old_0[12] , 
        \sr_new_0[12] , \sr_new_1[12] , \integral[6] , \integral[7] , 
        \integral[8] , \integral[9] , \integral[10] , \integral[11] , 
        \integral[12] , \integral[13] , \integral[14] , \integral[15] , 
        \integral[16] , \integral[17] , \integral[18] , \integral[19] , 
        \integral[20] , \integral[21] , \integral[22] , \integral[23] , 
        \integral[24] , \integral[25] , \integral_i[24] , 
        \integral_i[25] , \integral_0[25] , \integral_1[25] , 
        \derivative[12] , \sum[39] , \sum[14] , \sum[20] , \sum[19] , 
        \sum[22] , \sum[13] , \sum[17] , \sum[18] , \sum[21] , 
        \sum[23] , \sum[16] , \sum[15] , \sum[12] , \sum[11] , 
        \sum[6] , \sum[10] , \sum[9] , \sum[5] , \sum[8] , \sum[7] , 
        \sum[4] , \sum[2] , \sum[1] , \sum[0] , \sum[3] , \sum_0[39] , 
        \sum_1[39] , \sum_2[39] , vd_done, \off_div[0] , \off_div[1] , 
        \off_div[2] , \off_div[3] , \off_div[4] , \off_div[5] , 
        \off_div[6] , \off_div[7] , \off_div[8] , \off_div[9] , 
        \off_div[10] , \off_div[11] , \off_div[12] , \off_div[13] , 
        \off_div[14] , \off_div[15] , \off_div[16] , \off_div[17] , 
        \off_div[18] , \off_div[19] , \off_div[20] , \off_div[21] , 
        \off_div[22] , \off_div[23] , \off_div[24] , \off_div[25] , 
        \off_div[26] , \off_div[27] , \off_div[28] , \off_div[29] , 
        \off_div[30] , \off_div[31] , GND, VCC;
    
    pwm_ctl_400s_32s_13s_0_1_2_3 PWM_CTL (.sum_8(\sum[8] ), .sum_39(
        \sum[39] ), .sum_9(\sum[9] ), .sum_10(\sum[10] ), .sum_11(
        \sum[11] ), .sum_12(\sum[12] ), .sum_13(\sum[13] ), .sum_14(
        \sum[14] ), .sum_16(\sum[16] ), .sum_18(\sum[18] ), .sum_19(
        \sum[19] ), .sum_20(\sum[20] ), .sum_21(\sum[21] ), .sum_23(
        \sum[23] ), .sum_22(\sum[22] ), .sum_17(\sum[17] ), .sum_15(
        \sum[15] ), .sum_1_d0(\sum[1] ), .sum_0_d0(\sum[0] ), 
        .sum_2_d0(\sum[2] ), .sum_7(\sum[7] ), .sum_6(\sum[6] ), 
        .sum_4(\sum[4] ), .sum_3(\sum[3] ), .sum_5(\sum[5] ), .off_div({
        \off_div[31] , \off_div[30] , \off_div[29] , \off_div[28] , 
        \off_div[27] , \off_div[26] , \off_div[25] , \off_div[24] , 
        \off_div[23] , \off_div[22] , \off_div[21] , \off_div[20] , 
        \off_div[19] , \off_div[18] , \off_div[17] , \off_div[16] , 
        \off_div[15] , \off_div[14] , \off_div[13] , \off_div[12] , 
        \off_div[11] , \off_div[10] , \off_div[9] , \off_div[8] , 
        \off_div[7] , \off_div[6] , \off_div[5] , \off_div[4] , 
        \off_div[3] , \off_div[2] , \off_div[1] , \off_div[0] }), 
        .sum_2_0(\sum_2[39] ), .sum_1_0(\sum_1[39] ), .sum_0_0(
        \sum_0[39] ), .state({\state[1] , \state[0] }), .n_rst_c(
        n_rst_c), .clk_c(clk_c), .pwm_enable(pwm_enable));
    integral_calc_13s_4_1 AVG_CALC (.avg_old({\avg_old[11] , 
        \avg_old[10] , \avg_old[9] , \avg_old[8] , \avg_old[7] , 
        \avg_old[6] , \avg_old[5] , \avg_old[4] , \avg_old[3] , 
        \avg_old[2] , \avg_old[1] , \avg_old[0] }), .avg_new({
        \avg_new[11] , \avg_new[10] , \avg_new[9] , \avg_new[8] , 
        \avg_new[7] , \avg_new[6] , \avg_new[5] , \avg_new[4] , 
        \avg_new[3] , \avg_new[2] , \avg_new[1] , \avg_new[0] }), 
        .LED_33_0(LED_33_0), .choose({choose[2], choose[1], choose[0]})
        , .LED_5_0(LED_5_0), .LED_c_0(LED_c_0), .choose_0_0(choose_0_0)
        , .LED_15_0(LED_15_0), .LED_12_0(LED_12_0), .average({
        \average[6] , \average[5] , \average[4] , \average[3] , 
        \average[2] }), .LED_FB({LED_FB[7], LED_FB[6], LED_FB[5], 
        \LED_FB[4] , LED_FB[3], LED_FB[2], LED_FB[1], LED_FB[0]}), 
        .LED_FB_i_0(\LED_FB_i[5] ), .calc_avg(calc_avg), .avg_done(
        avg_done), .n_rst_c(n_rst_c), .clk_c(clk_c));
    error_sr_13s_5s_1 AVGSR (.cur_vd({\cur_vd[11] , \cur_vd[10] , 
        \cur_vd[9] , \cur_vd[8] , \cur_vd[7] , \cur_vd[6] , 
        \cur_vd[5] , \cur_vd[4] , \cur_vd[3] , \cur_vd[2] , 
        \cur_vd[1] , \cur_vd[0] }), .avg_new({\avg_new[11] , 
        \avg_new[10] , \avg_new[9] , \avg_new[8] , \avg_new[7] , 
        \avg_new[6] , \avg_new[5] , \avg_new[4] , \avg_new[3] , 
        \avg_new[2] , \avg_new[1] , \avg_new[0] }), .avg_old({
        \avg_old[11] , \avg_old[10] , \avg_old[9] , \avg_old[8] , 
        \avg_old[7] , \avg_old[6] , \avg_old[5] , \avg_old[4] , 
        \avg_old[3] , \avg_old[2] , \avg_old[1] , \avg_old[0] }), 
        .avg_enable(avg_enable), .avg_enable_1(avg_enable_1), 
        .avg_enable_0(avg_enable_0), .n_rst_c(n_rst_c), .clk_c(clk_c));
    error_sr_13s_64s_1 INTSR (.sr_old({\sr_old[12] , \sr_old[11] , 
        \sr_old[10] , \sr_old[9] , \sr_old[8] , \sr_old[7] , 
        \sr_old[6] , \sr_old[5] , \sr_old[4] , \sr_old[3] , 
        \sr_old[2] , \sr_old[1] , \sr_old[0] }), .sr_new({\sr_new[12] , 
        \sr_new[11] , \sr_new[10] , \sr_new[9] , \sr_new[8] , 
        \sr_new[7] , \sr_new[6] , \sr_new[5] , \sr_new[4] , 
        \sr_new[3] , \sr_new[2] , \sr_new[1] , \sr_new[0] }), 
        .cur_error({\cur_error[12] , \cur_error[11] , \cur_error[10] , 
        \cur_error[9] , \cur_error[8] , \cur_error[7] , \cur_error[6] , 
        \cur_error[5] , \cur_error[4] , \cur_error[3] , \cur_error[2] , 
        \cur_error[1] , \cur_error[0] }), .sr_prev({\sr_prev[12] , 
        \sr_prev[11] , \sr_prev[10] , \sr_prev[9] , \sr_prev[8] , 
        \sr_prev[7] , \sr_prev[6] , \sr_prev[5] , \sr_prev[4] , 
        \sr_prev[3] , \sr_prev[2] , \sr_prev[1] , \sr_prev[0] }), 
        .sr_old_0_0(\sr_old_0[12] ), .sr_new_0_0(\sr_new_0[12] ), 
        .sr_new_1_0(\sr_new_1[12] ), .int_enable_11(int_enable_11), 
        .int_enable_29(int_enable_29), .int_enable_19(int_enable_19), 
        .int_enable_8(int_enable_8), .int_enable_4(int_enable_4), 
        .int_enable_28(int_enable_28), .int_enable_17(int_enable_17), 
        .int_enable_26(int_enable_26), .int_enable_9(int_enable_9), 
        .int_enable_18(int_enable_18), .int_enable_21(int_enable_21), 
        .int_enable_20(int_enable_20), .int_enable_27(int_enable_27), 
        .int_enable_31(int_enable_31), .int_enable_30(int_enable_30), 
        .int_enable_5(int_enable_5), .int_enable_3(int_enable_3), 
        .int_enable_2(int_enable_2), .int_enable_14(int_enable_14), 
        .int_enable_13(int_enable_13), .int_enable_23(int_enable_23), 
        .int_enable_12(int_enable_12), .int_enable_32(int_enable_32), 
        .int_enable_1(int_enable_1), .int_enable_7(int_enable_7), 
        .int_enable_6(int_enable_6), .int_enable_22(int_enable_22), 
        .int_enable_16(int_enable_16), .int_enable_15(int_enable_15), 
        .int_enable_10(int_enable_10), .int_enable_25(int_enable_25), 
        .int_enable_24(int_enable_24), .int_enable_33(int_enable_33), 
        .int_enable(int_enable), .int_enable_0(int_enable_0), .n_rst_c(
        n_rst_c), .clk_c(clk_c));
    controller_Z1_4_1 CONTROLLER (.state_0_d0(\state[1] ), .state_0_0(
        \state[0] ), .pwm_chg(pwm_chg), .int_done(int_done), .sig_prev(
        sig_prev), .sig_old_i_0(sig_old_i_0), .avg_done(avg_done), 
        .int_enable(int_enable), .vd_rdy(vd_rdy), .sum_rdy(sum_rdy), 
        .deriv_enable(deriv_enable), .calc_avg(calc_avg), .calc_int(
        calc_int), .pwm_enable(pwm_enable), .sum_enable(sum_enable), 
        .avg_enable(avg_enable), .pwm_chg_0(pwm_chg_0), .int_enable_0(
        int_enable_0), .int_enable_1(int_enable_1), .int_enable_2(
        int_enable_2), .int_enable_3(int_enable_3), .int_enable_4(
        int_enable_4), .int_enable_5(int_enable_5), .int_enable_6(
        int_enable_6), .int_enable_7(int_enable_7), .int_enable_8(
        int_enable_8), .int_enable_9(int_enable_9), .int_enable_10(
        int_enable_10), .int_enable_11(int_enable_11), .int_enable_12(
        int_enable_12), .int_enable_13(int_enable_13), .int_enable_14(
        int_enable_14), .int_enable_15(int_enable_15), .int_enable_16(
        int_enable_16), .int_enable_17(int_enable_17), .int_enable_18(
        int_enable_18), .int_enable_19(int_enable_19), .int_enable_20(
        int_enable_20), .int_enable_21(int_enable_21), .int_enable_22(
        int_enable_22), .int_enable_23(int_enable_23), .int_enable_24(
        int_enable_24), .int_enable_25(int_enable_25), .int_enable_26(
        int_enable_26), .int_enable_27(int_enable_27), .int_enable_28(
        int_enable_28), .int_enable_29(int_enable_29), .int_enable_30(
        int_enable_30), .int_enable_31(int_enable_31), .int_enable_32(
        int_enable_32), .int_enable_33(int_enable_33), .avg_enable_0(
        avg_enable_0), .n_rst_c(n_rst_c), .clk_c(clk_c), .avg_enable_1(
        avg_enable_1), .calc_error(calc_error));
    sig_gen_4 FM_CYCLE (.primary_fb_c(primary_fb_c), .n_rst_c(n_rst_c), 
        .clk_c(clk_c), .sig_old_i_0(sig_old_i_0), .sig_prev(sig_prev));
    pid_sum_13s_4_1 SUM (.integral_i({\integral_i[25] , 
        \integral_i[24] }), .integral({\integral[25] , \integral[24] , 
        \integral[23] , \integral[22] , \integral[21] , \integral[20] , 
        \integral[19] , \integral[18] , \integral[17] , \integral[16] , 
        \integral[15] , \integral[14] , \integral[13] , \integral[12] , 
        \integral[11] , \integral[10] , \integral[9] , \integral[8] , 
        \integral[7] , \integral[6] }), .sr_new({\sr_new[12] , 
        \sr_new[11] , \sr_new[10] , \sr_new[9] , \sr_new[8] , 
        \sr_new[7] , \sr_new[6] , \sr_new[5] , \sr_new[4] , 
        \sr_new[3] , \sr_new[2] , \sr_new[1] , \sr_new[0] }), 
        .derivative_0(\derivative[12] ), .sr_new_1_0(\sr_new_1[12] ), 
        .sr_new_0_0(\sr_new_0[12] ), .integral_1_0(\integral_1[25] ), 
        .integral_0_0(\integral_0[25] ), .sum_39(\sum[39] ), .sum_14(
        \sum[14] ), .sum_20(\sum[20] ), .sum_19(\sum[19] ), .sum_22(
        \sum[22] ), .sum_13(\sum[13] ), .sum_17(\sum[17] ), .sum_18(
        \sum[18] ), .sum_21(\sum[21] ), .sum_23(\sum[23] ), .sum_16(
        \sum[16] ), .sum_15(\sum[15] ), .sum_12(\sum[12] ), .sum_11(
        \sum[11] ), .sum_6(\sum[6] ), .sum_10(\sum[10] ), .sum_9(
        \sum[9] ), .sum_5(\sum[5] ), .sum_8(\sum[8] ), .sum_7(\sum[7] )
        , .sum_4(\sum[4] ), .sum_2_d0(\sum[2] ), .sum_1_d0(\sum[1] ), 
        .sum_0_d0(\sum[0] ), .sum_3(\sum[3] ), .sum_0_0(\sum_0[39] ), 
        .sum_1_0(\sum_1[39] ), .sum_2_0(\sum_2[39] ), .sum_enable(
        sum_enable), .sum_rdy(sum_rdy), .n_rst_c(n_rst_c), .clk_c(
        clk_c));
    sig_gen_3 VD_SIG (.vd_done(vd_done), .n_rst_c(n_rst_c), .clk_c(
        clk_c), .vd_rdy(vd_rdy));
    spi_rx_12s_3_0 SPI (.cur_vd({\cur_vd[11] , \cur_vd[10] , 
        \cur_vd[9] , \cur_vd[8] , \cur_vd[7] , \cur_vd[6] , 
        \cur_vd[5] , \cur_vd[4] , \cur_vd[3] , \cur_vd[2] , 
        \cur_vd[1] , \cur_vd[0] }), .vd_done(vd_done), .cs_i_1_i(
        cs_i_1_i), .sck_33_c(sck_33_c), .n_rst_c(n_rst_c), .din_fb_c(
        din_fb_c));
    integral_calc_13s_0_4_1 INTCALC (.sr_old({\sr_old[12] , 
        \sr_old[11] , \sr_old[10] , \sr_old[9] , \sr_old[8] , 
        \sr_old[7] , \sr_old[6] , \sr_old[5] , \sr_old[4] , 
        \sr_old[3] , \sr_old[2] , \sr_old[1] , \sr_old[0] }), .sr_new({
        \sr_new[12] , \sr_new[11] , \sr_new[10] , \sr_new[9] , 
        \sr_new[8] , \sr_new[7] , \sr_new[6] , \sr_new[5] , 
        \sr_new[4] , \sr_new[3] , \sr_new[2] , \sr_new[1] , 
        \sr_new[0] }), .sr_new_0_0(\sr_new_0[12] ), .sr_new_1_0(
        \sr_new_1[12] ), .integral({\integral[25] , \integral[24] , 
        \integral[23] , \integral[22] , \integral[21] , \integral[20] , 
        \integral[19] , \integral[18] , \integral[17] , \integral[16] , 
        \integral[15] , \integral[14] , \integral[13] , \integral[12] , 
        \integral[11] , \integral[10] , \integral[9] , \integral[8] , 
        \integral[7] , \integral[6] }), .sr_old_0_0(\sr_old_0[12] ), 
        .integral_i({\integral_i[25] , \integral_i[24] }), 
        .integral_0_0(\integral_0[25] ), .integral_1_0(
        \integral_1[25] ), .calc_int(calc_int), .int_done(int_done), 
        .n_rst_c(n_rst_c), .clk_c(clk_c));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    error_calc_13s_12s_4_1 EC (.cur_error({\cur_error[12] , 
        \cur_error[11] , \cur_error[10] , \cur_error[9] , 
        \cur_error[8] , \cur_error[7] , \cur_error[6] , \cur_error[5] , 
        \cur_error[4] , \cur_error[3] , \cur_error[2] , \cur_error[1] , 
        \cur_error[0] }), .LED_FB_i_0(\LED_FB_i[5] ), .LED_FB({
        LED_FB[7], LED_FB[6], LED_FB[5], \LED_FB[4] , LED_FB[3], 
        LED_FB[2], LED_FB[1], LED_FB[0]}), .average({\average[6] , 
        \average[5] , \average[4] , \average[3] , \average[2] }), 
        .calc_error(calc_error), .n_rst_c(n_rst_c), .clk_c(clk_c));
    derivative_calc_13s_4_1 DCALC (.derivative_0(\derivative[12] ), 
        .sr_new({\sr_new[12] , \sr_new[11] , \sr_new[10] , \sr_new[9] , 
        \sr_new[8] , \sr_new[7] , \sr_new[6] , \sr_new[5] , 
        \sr_new[4] , \sr_new[3] , \sr_new[2] , \sr_new[1] , 
        \sr_new[0] }), .sr_prev({\sr_prev[12] , \sr_prev[11] , 
        \sr_prev[10] , \sr_prev[9] , \sr_prev[8] , \sr_prev[7] , 
        \sr_prev[6] , \sr_prev[5] , \sr_prev[4] , \sr_prev[3] , 
        \sr_prev[2] , \sr_prev[1] , \sr_prev[0] }), .deriv_enable(
        deriv_enable), .n_rst_c(n_rst_c), .clk_c(clk_c));
    pwm_tx_400s_32s_13s_10_1000000s_45s_1_0 PWM_TX (.off_div({
        \off_div[31] , \off_div[30] , \off_div[29] , \off_div[28] , 
        \off_div[27] , \off_div[26] , \off_div[25] , \off_div[24] , 
        \off_div[23] , \off_div[22] , \off_div[21] , \off_div[20] , 
        \off_div[19] , \off_div[18] , \off_div[17] , \off_div[16] , 
        \off_div[15] , \off_div[14] , \off_div[13] , \off_div[12] , 
        \off_div[11] , \off_div[10] , \off_div[9] , \off_div[8] , 
        \off_div[7] , \off_div[6] , \off_div[5] , \off_div[4] , 
        \off_div[3] , \off_div[2] , \off_div[1] , \off_div[0] }), 
        .act_ctl_5_i(act_ctl_5_i), .act_ctl_5_3(act_ctl_5_3), 
        .act_ctl_5_0(act_ctl_5_0), .pwm_chg_0(pwm_chg_0), .pwm_chg(
        pwm_chg), .n_rst_c(n_rst_c), .clk_c(clk_c), .act_ctl_5_2(
        act_ctl_5_2), .act_ctl_5_1(act_ctl_5_1), .act_ctl_5_9(
        act_ctl_5_9), .act_ctl_5_8(act_ctl_5_8), .act_ctl_5(act_ctl_5), 
        .primary_fb_c(primary_fb_c));
    spi_clk_11s_3_0 SPICLK (.sck_33_c(sck_33_c), .n_rst_c(n_rst_c), 
        .clk_c(clk_c));
    
endmodule


module PSU_controller(
       act_ctl_5,
       act_ctl_5_i,
       act_ctl_5_0,
       act_ctl_5_1,
       act_ctl_5_2,
       act_ctl_5_3,
       act_ctl_5_4,
       act_ctl_5_5,
       act_ctl_5_6,
       act_ctl_5_7,
       act_ctl_5_8,
       n_rst_c,
       clk_c,
       act_ctl_5_9
    );
output act_ctl_5;
output act_ctl_5_i;
output act_ctl_5_0;
output act_ctl_5_1;
output act_ctl_5_2;
output act_ctl_5_3;
output act_ctl_5_4;
output act_ctl_5_5;
output act_ctl_5_6;
output act_ctl_5_7;
output act_ctl_5_8;
input  n_rst_c;
input  clk_c;
output act_ctl_5_9;

    wire N_7, cnt_e11_0_0, \cnt[10]_net_1 , \cnt[11]_net_1 , N_66, 
        N_68, cnt_e10_0_a3_0_0, N_36, cnt_e11_0_a3_1_0, N_69, 
        \cnt[9]_net_1 , N_35, N_76, N_71, N_116, cnt_e9, N_70, cnt_e11, 
        N_109, N_27, \cnt[0]_net_1 , \cnt_i_0[1] , N_28, \cnt_i_0[2] , 
        N_29, \cnt_i_0[3] , N_30, \cnt_i_0[4] , N_31, \cnt[5]_net_1 , 
        N_32, \cnt[6]_net_1 , \cnt[7]_net_1 , \cnt[8]_net_1 , cnt_e10, 
        cnt_e8_0_a3_1_0, cnt_e8_0_a3_0, cnt_e1_i_0, cnt_e2_i_0, 
        cnt_e3_i_0, cnt_e6_i_0, cnt_e4_i_0, cnt_e5_i_0, 
        un1_cntlto11_i_a2_2, un1_cntlto11_i_a2_1, un1_cntlto11_i_a2_0, 
        cnt_e8, N_72, N_73, N_74, N_13, N_75, N_122, N_78, N_15, N_17, 
        N_19, N_21, N_23, N_25, \state_ns[1] , \state[1]_net_1 , 
        cnt_e0, GND, VCC;
    
    OR3 \cnt_RNO[8]  (.A(N_72), .B(N_73), .C(N_74), .Y(cnt_e8));
    NOR3C \cnt_RNIP7131[5]  (.A(un1_cntlto11_i_a2_1), .B(
        un1_cntlto11_i_a2_0), .C(un1_cntlto11_i_a2_2), .Y(N_76));
    DFN1C0 \state_7[0]  (.D(N_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        act_ctl_5_7));
    DFN1C0 \state_3[0]  (.D(N_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        act_ctl_5_3));
    AX1 \cnt_RNO_0[3]  (.A(N_28), .B(act_ctl_5_1), .C(\cnt_i_0[3] ), 
        .Y(cnt_e3_i_0));
    OR3B \cnt_RNI1KKG[8]  (.A(\cnt[7]_net_1 ), .B(\cnt[8]_net_1 ), .C(
        N_32), .Y(N_35));
    OR2 \cnt_RNO[2]  (.A(cnt_e2_i_0), .B(N_122), .Y(N_23));
    DFN1P0 \cnt[2]  (.D(N_23), .CLK(clk_c), .PRE(n_rst_c), .Q(
        \cnt_i_0[2] ));
    DFN1C0 \cnt[8]  (.D(cnt_e8), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \cnt[8]_net_1 ));
    DFN1P0 \cnt[1]  (.D(N_25), .CLK(clk_c), .PRE(n_rst_c), .Q(
        \cnt_i_0[1] ));
    AX1 \cnt_RNO_0[4]  (.A(N_29), .B(act_ctl_5_0), .C(\cnt_i_0[4] ), 
        .Y(cnt_e4_i_0));
    DFN1C0 \cnt[11]  (.D(cnt_e11), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \cnt[11]_net_1 ));
    AX1A \cnt_RNO_0[6]  (.A(N_31), .B(act_ctl_5_1), .C(\cnt[6]_net_1 ), 
        .Y(cnt_e6_i_0));
    OR2 \cnt_RNIJI79[4]  (.A(\cnt_i_0[4] ), .B(N_29), .Y(N_30));
    NOR3B \cnt_RNO_2[8]  (.A(\cnt[7]_net_1 ), .B(cnt_e8_0_a3_1_0), .C(
        N_32), .Y(N_74));
    NOR3B \cnt_RNO_1[7]  (.A(\cnt[7]_net_1 ), .B(act_ctl_5_1), .C(N_32)
        , .Y(N_78));
    OR2 \cnt_RNO[3]  (.A(cnt_e3_i_0), .B(N_122), .Y(N_21));
    NOR2A \cnt_RNO_1[8]  (.A(\cnt[8]_net_1 ), .B(act_ctl_5_4), .Y(N_73)
        );
    NOR2B \cnt_RNI3NNE[11]  (.A(\cnt[11]_net_1 ), .B(\cnt[7]_net_1 ), 
        .Y(un1_cntlto11_i_a2_0));
    VCC VCC_i (.Y(VCC));
    OR2 \cnt_RNO[1]  (.A(cnt_e1_i_0), .B(N_122), .Y(N_25));
    NOR2A \cnt_RNO_3[8]  (.A(\cnt[8]_net_1 ), .B(N_76), .Y(
        cnt_e8_0_a3_0));
    DFN1C0 \cnt[6]  (.D(N_15), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \cnt[6]_net_1 ));
    DFN1C0 \state_0[0]  (.D(N_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        act_ctl_5_0));
    DFN1P0 \cnt[4]  (.D(N_19), .CLK(clk_c), .PRE(n_rst_c), .Q(
        \cnt_i_0[4] ));
    DFN1C0 \state_2[0]  (.D(N_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        act_ctl_5_2));
    DFN1C0 \cnt[9]  (.D(cnt_e9), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \cnt[9]_net_1 ));
    DFN1C0 \state_4[0]  (.D(N_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        act_ctl_5_4));
    AXOI4 \cnt_RNO[0]  (.A(N_76), .B(act_ctl_5_0), .C(\cnt[0]_net_1 ), 
        .Y(cnt_e0));
    DFN1C0 \cnt[0]  (.D(cnt_e0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \cnt[0]_net_1 ));
    DFN1C0 \state_6[0]  (.D(N_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        act_ctl_5_6));
    AO1C \state_0_RNIOV4M1[0]  (.A(N_76), .B(N_36), .C(act_ctl_5_0), 
        .Y(N_109));
    OR2 \cnt_RNO[4]  (.A(cnt_e4_i_0), .B(N_122), .Y(N_19));
    OA1 \cnt_RNIIOH5[5]  (.A(\cnt[5]_net_1 ), .B(\cnt[6]_net_1 ), .C(
        \cnt[8]_net_1 ), .Y(un1_cntlto11_i_a2_2));
    NOR2B \cnt_RNI4ONE[9]  (.A(\cnt[10]_net_1 ), .B(\cnt[9]_net_1 ), 
        .Y(un1_cntlto11_i_a2_1));
    DFN1C0 \state[0]  (.D(N_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        act_ctl_5));
    NOR2 \cnt_RNO[6]  (.A(cnt_e6_i_0), .B(N_122), .Y(N_15));
    OA1C \cnt_RNO_0[7]  (.A(act_ctl_5_0), .B(N_32), .C(\cnt[7]_net_1 ), 
        .Y(N_75));
    OR3 \cnt_RNO[9]  (.A(N_69), .B(N_70), .C(N_71), .Y(cnt_e9));
    INV \state_RNIHMTD[0]  (.A(act_ctl_5), .Y(act_ctl_5_i));
    GND GND_i (.Y(GND));
    NOR2B \state_4_RNITC181[0]  (.A(N_76), .B(act_ctl_5_4), .Y(N_122));
    OR2A \cnt_RNI81UC[6]  (.A(\cnt[6]_net_1 ), .B(N_31), .Y(N_32));
    NOR2A \state_4_RNITC181_0[0]  (.A(act_ctl_5_4), .B(N_76), .Y(N_116)
        );
    NOR3A \cnt_RNO_2[9]  (.A(N_116), .B(\cnt[9]_net_1 ), .C(N_35), .Y(
        N_71));
    NOR3B \cnt_RNO_0[9]  (.A(\cnt[9]_net_1 ), .B(N_35), .C(N_76), .Y(
        N_69));
    DFN1C0 \cnt[7]  (.D(N_13), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \cnt[7]_net_1 ));
    DFN1C0 \cnt[10]  (.D(cnt_e10), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \cnt[10]_net_1 ));
    AX1C \cnt_RNO_0[1]  (.A(\cnt[0]_net_1 ), .B(act_ctl_5_0), .C(
        \cnt_i_0[1] ), .Y(cnt_e1_i_0));
    NOR2A \cnt_RNO_1[11]  (.A(cnt_e11_0_a3_1_0), .B(N_36), .Y(N_66));
    NOR2 \cnt_RNO[5]  (.A(cnt_e5_i_0), .B(N_122), .Y(N_17));
    OR2 \cnt_RNI28H5[2]  (.A(\cnt_i_0[2] ), .B(N_27), .Y(N_28));
    DFN1C0 \state[1]  (.D(\state_ns[1] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[1]_net_1 ));
    OA1A \cnt_RNO_0[8]  (.A(\cnt[7]_net_1 ), .B(N_32), .C(
        cnt_e8_0_a3_0), .Y(N_72));
    DFN1P0 \cnt[3]  (.D(N_21), .CLK(clk_c), .PRE(n_rst_c), .Q(
        \cnt_i_0[3] ));
    NOR2B \cnt_RNO_2[11]  (.A(\cnt[10]_net_1 ), .B(N_116), .Y(
        cnt_e11_0_a3_1_0));
    NOR2 \state_RNIF4VL1[1]  (.A(\state[1]_net_1 ), .B(N_122), .Y(N_7));
    DFN1C0 \state_9[0]  (.D(N_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        act_ctl_5_9));
    NOR2A \cnt_RNO_1[10]  (.A(N_116), .B(\cnt[10]_net_1 ), .Y(
        cnt_e10_0_a3_0_0));
    AO1A \cnt_RNO_0[11]  (.A(\cnt[10]_net_1 ), .B(\cnt[11]_net_1 ), .C(
        N_66), .Y(cnt_e11_0_0));
    DFN1C0 \state_1[0]  (.D(N_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        act_ctl_5_1));
    AO1 \cnt_RNO[11]  (.A(N_109), .B(\cnt[11]_net_1 ), .C(cnt_e11_0_0), 
        .Y(cnt_e11));
    NOR2A \cnt_RNO_1[9]  (.A(\cnt[9]_net_1 ), .B(act_ctl_5_6), .Y(N_70)
        );
    AX1 \cnt_RNO_0[2]  (.A(N_27), .B(act_ctl_5_0), .C(\cnt_i_0[2] ), 
        .Y(cnt_e2_i_0));
    AO1 \cnt_RNO[10]  (.A(N_109), .B(\cnt[10]_net_1 ), .C(N_68), .Y(
        cnt_e10));
    AX1A \cnt_RNO_0[5]  (.A(N_30), .B(act_ctl_5_0), .C(\cnt[5]_net_1 ), 
        .Y(cnt_e5_i_0));
    OR2A \cnt_RNIB4M3[1]  (.A(\cnt[0]_net_1 ), .B(\cnt_i_0[1] ), .Y(
        N_27));
    OR2A \cnt_RNIDP2B[5]  (.A(\cnt[5]_net_1 ), .B(N_30), .Y(N_31));
    NOR2A \cnt_RNO_0[10]  (.A(cnt_e10_0_a3_0_0), .B(N_36), .Y(N_68));
    DFN1C0 \cnt[5]  (.D(N_17), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \cnt[5]_net_1 ));
    DFN1C0 \state_8[0]  (.D(N_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        act_ctl_5_8));
    DFN1C0 \state_5[0]  (.D(N_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        act_ctl_5_5));
    OR2 \cnt_RNIQCC7[3]  (.A(\cnt_i_0[3] ), .B(N_28), .Y(N_29));
    AXOI5 \state_RNO[1]  (.A(N_76), .B(act_ctl_5_0), .C(
        \state[1]_net_1 ), .Y(\state_ns[1] ));
    NOR2A \cnt_RNO_4[8]  (.A(N_116), .B(\cnt[8]_net_1 ), .Y(
        cnt_e8_0_a3_1_0));
    OR2A \cnt_RNIVUFI[9]  (.A(\cnt[9]_net_1 ), .B(N_35), .Y(N_36));
    NOR3 \cnt_RNO[7]  (.A(N_75), .B(N_122), .C(N_78), .Y(N_13));
    
endmodule


module pwm_ctl_400s_32s_13s_0_1_2_2(
       sum_8,
       sum_39,
       sum_12,
       sum_14,
       sum_9,
       sum_10,
       sum_11,
       sum_13,
       sum_15,
       sum_18,
       sum_21,
       sum_22,
       sum_23,
       sum_16,
       sum_17,
       sum_20,
       sum_19,
       sum_1_d0,
       sum_0_d0,
       sum_2_d0,
       sum_7,
       sum_6,
       sum_5,
       sum_4,
       sum_3,
       off_div,
       sum_2_0,
       sum_1_0,
       sum_0_0,
       n_rst_c,
       clk_c,
       pwm_rdy,
       pwm_enable
    );
input  sum_8;
input  sum_39;
input  sum_12;
input  sum_14;
input  sum_9;
input  sum_10;
input  sum_11;
input  sum_13;
input  sum_15;
input  sum_18;
input  sum_21;
input  sum_22;
input  sum_23;
input  sum_16;
input  sum_17;
input  sum_20;
input  sum_19;
input  sum_1_d0;
input  sum_0_d0;
input  sum_2_d0;
input  sum_7;
input  sum_6;
input  sum_5;
input  sum_4;
input  sum_3;
output [31:0] off_div;
input  sum_2_0;
input  sum_1_0;
input  sum_0_0;
input  n_rst_c;
input  clk_c;
output pwm_rdy;
input  pwm_enable;

    wire \state_d_0[2] , \state[1]_net_1 , \state[0]_net_1 , 
        un1_state_2_0, un5lt31, next_off_div_2_sqmuxa_11, N_16, 
        \DWACT_FINC_E[4] , N_13, \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , 
        ADD_32x32_fast_I321_Y_0, ADD_32x32_fast_I258_Y_3, N610, N625, 
        ADD_32x32_fast_I258_Y_2, N482, ADD_32x32_fast_I258_Y_0, N551, 
        ADD_32x32_fast_I320_Y_0, ADD_32x32_fast_I313_Y_0, 
        ADD_32x32_fast_I259_Y_3, N612, N627, ADD_32x32_fast_I259_Y_2, 
        N484, ADD_32x32_fast_I259_Y_0, N553, 
        ADD_32x32_fast_I258_un1_Y_0, N626, ADD_32x32_fast_I319_Y_0, 
        ADD_32x32_fast_I318_Y_0, ADD_32x32_fast_I317_Y_0, 
        ADD_32x32_fast_I316_Y_0, ADD_32x32_fast_I315_Y_0, 
        ADD_32x32_fast_I314_Y_0, ADD_32x32_fast_I266_Y_0, N641, 
        ADD_32x32_fast_I260_Y_2, N614, N629, ADD_32x32_fast_I260_Y_1, 
        N486, N555, ADD_32x32_fast_I261_Y_2, N616, N631, 
        ADD_32x32_fast_I261_Y_1, N488, N557, ADD_32x32_fast_I312_Y_0, 
        ADD_32x32_fast_I304_Y_0, \sum_adj[22]_net_1 , 
        ADD_32x32_fast_I259_un1_Y_0, N628, ADD_32x32_fast_I262_Y_1, 
        N618, N633, ADD_32x32_fast_I262_Y_0, N559, 
        ADD_32x32_fast_I310_Y_0, ADD_32x32_fast_I311_Y_0, 
        ADD_32x32_fast_I309_Y_0, ADD_32x32_fast_I266_un1_Y_0, N642, 
        ADD_32x32_fast_I264_Y_1, N622, N637, ADD_32x32_fast_I264_Y_0, 
        N563, ADD_32x32_fast_I263_Y_1, N620, N635, 
        ADD_32x32_fast_I263_Y_0, N561, ADD_32x32_fast_I265_Y_0, N565, 
        ADD_32x32_fast_I306_Y_0, ADD_32x32_fast_I307_Y_0, 
        ADD_32x32_fast_I308_Y_0, ADD_32x32_fast_I303_Y_0, 
        \un1_sum_adj[13] , ADD_32x32_fast_I302_Y_0, \un1_sum_adj[12] , 
        ADD_32x32_fast_I260_un1_Y_0, N630, ADD_32x32_fast_I261_un1_Y_0, 
        N632, ADD_32x32_fast_I301_Y_0, \un1_sum_adj[11] , 
        ADD_32x32_fast_I262_un1_Y_0, N634, ADD_32x32_fast_I269_Y_0, 
        N647, ADD_32x32_fast_I270_Y_0, N649, ADD_32x32_fast_I299_Y_0, 
        \un1_sum_adj[9] , ADD_32x32_fast_I300_Y_0, \un1_sum_adj[10] , 
        ADD_32x32_fast_I298_Y_0, \un1_sum_adj[8] , 
        ADD_32x32_fast_I265_un1_Y_0, N624, N640, 
        ADD_32x32_fast_I264_un1_Y_0, N638, ADD_32x32_fast_I263_un1_Y_0, 
        N636, ADD_32x32_fast_I296_Y_0, \un1_sum_adj[6] , 
        ADD_32x32_fast_I273_Y_0, ADD_32x32_fast_I273_un1_Y_0, N639, 
        ADD_32x32_fast_I272_Y_0, ADD_32x32_fast_I272_un1_Y_0, 
        ADD_32x32_fast_I271_Y_0, ADD_32x32_fast_I271_un1_Y_0, 
        ADD_32x32_fast_I294_Y_0, \un1_sum_adj[4] , 
        ADD_32x32_fast_I295_Y_0, \un1_sum_adj[5] , 
        ADD_32x32_fast_I293_Y_0, \sum_adj[11]_net_1 , N590, N598, 
        \un1_sum_adj[0] , N538, N654, N586, N594, N601, 
        ADD_32x32_fast_I292_Y_0, \sum_adj[10]_net_1 , 
        next_off_div_2_sqmuxa_10, next_off_div37, 
        next_off_div_2_sqmuxa_7, next_off_div_2_sqmuxa_6, 
        next_off_div_2_sqmuxa_8, un1_off_divlto31_10, 
        next_off_div_2_sqmuxa_5, next_off_div_2_sqmuxa_2, 
        un1_off_divlto31_9, next_off_div_2_sqmuxa_1, 
        ADD_32x32_fast_I291_Y_0, \un1_sum_adj[1] , un5lto20_2, 
        un5lto20_1, ADD_32x32_fast_I159_Y_0, N483, N487, 
        ADD_32x32_fast_I157_Y_1, ADD_32x32_fast_I157_Y_0, N485, 
        ADD_32x32_fast_I155_Y_0, ADD_32x32_fast_I161_Y_0, N489, 
        un5lto14_2, un5lto14_1, un1_off_divlto31_22, 
        un1_off_divlto31_15, un1_off_divlto31_14, un1_off_divlto31_20, 
        un1_off_divlto31_21, un1_off_divlto31_13, un1_off_divlto31_12, 
        un1_off_divlto31_17, un1_off_divlt31, un1_off_divlto31_0, 
        un5lto9, un1_off_divlto31_8, un1_off_divlto31_6, 
        un1_off_divlto31_4, un1_off_divlto31_2, un5lto7_1, N495, N491, 
        I267_un1_Y, N644, N659, N767, I228_un1_Y, \un1_off_div_1[19] , 
        I270_un1_Y, N650, N599, N753, N787, N779, N655, 
        \un1_off_div_1[15] , \un1_sum_adj[15] , N781, N755, N790, N558, 
        \un1_off_div_1[18] , I236_un1_Y, N763, I224_un1_Y, I265_un1_Y, 
        N802, N749, N552, N751, N784, N493, N757, N793, N765, N657, 
        un5lt16, I269_un1_Y, N648, N663, \un1_off_div_1[20] , 
        \un1_off_div_1[17] , I238_un1_Y, un5lt9, un5lto4, un5lt4, 
        un1_off_div, \un1_off_div_1[0] , \un1_off_div_1[10] , N796, 
        \un1_off_div_1[7] , \un1_sum_adj[7] , \un1_off_div_1[5] , N661, 
        \un1_off_div_1[3] , N769, I230_un1_Y, I268_un1_Y, N646, N761, 
        N799, N759, \state_ns[0] , N_311_i, \nsum_adj_11[12] , I_35_0, 
        \nsum_adj_11[8] , I_23_2, \nsum_adj_11[14] , I_40_0, 
        \next_off_div[2] , \state_d[2] , \next_off_div[9] , 
        \next_off_div[11] , \next_off_div[12] , \next_off_div[13] , 
        \next_off_div[21] , \next_off_div[25] , \next_off_div[26] , 
        N383, N386, N387, N390, N392, N393, N398, N399, N404, N405, 
        N521, N411, N522, N523, N524, N401, N525, N526, N527, N528, 
        N395, N529, N531, N532, N389, N533, N534, N535, N536, N537, 
        \sum_adj[8]_net_1 , N580, N515, N519, N584, N587, N588, N589, 
        N592, N593, N596, N597, I150_un1_Y, N564, N572, N579, N571, 
        N645, N518, N514, N416, N417, N407, N413, N419, N422, N423, 
        N426, N516, N517, N581, N520, N582, N583, N585, N562, 
        I184_un1_Y, N574, N573, N653, \nsum_adj_11[9] , I_26_0, 
        \nsum_adj_11[10] , I_28_0, \nsum_adj_11[11] , I_32_0, 
        \nsum_adj_11[13] , I_37_0, \nsum_adj_11[15] , I_43_0, 
        \nsum_adj_11[18] , I_53_0, \nsum_adj_11[21] , I_62_0, 
        \nsum_adj_11[22] , I_65_0, \nsum_adj_11[23] , I_70_0, 
        \sum_adj[21]_net_1 , \sum_adj[20]_net_1 , \sum_adj[19]_net_1 , 
        \sum_adj[18]_net_1 , \sum_adj[16]_net_1 , \sum_adj[15]_net_1 , 
        \sum_adj[13]_net_1 , \sum_adj[9]_net_1 , \next_off_div[5] , 
        next_off_div_0_sqmuxa, \next_off_div[3] , \next_off_div[0] , 
        state_176_d, N566, N504, N500, N497, N501, N496, N492, 
        \next_off_div[7] , next_off_div_1_sqmuxa, \next_off_div[10] , 
        \next_off_div[17] , \next_off_div[20] , \nsum_adj_11[16] , 
        I_46_0, un1_state_2, un5lt14, \sum_adj[14]_net_1 , I247_un1_Y, 
        N651, N570, N569, \next_off_div[6] , \next_off_div[27] , 
        \next_off_div[23] , N560, \next_off_div[30] , 
        \next_off_div[31] , \sum_adj[17]_net_1 , N591, N576, N575, 
        N568, N567, N511, N510, N503, N507, N506, N502, N410, 
        \next_off_div[24] , N428, N432, N505, N509, N577, N578, 
        \next_off_div[18] , \next_off_div[28] , N429, N508, N425, 
        \sum_adj[23]_net_1 , \next_off_div[15] , I249_un1_Y, N513, 
        N512, \next_off_div[29] , \next_off_div[16] , 
        \next_off_div[14] , \next_off_div[8] , \next_off_div[1] , N490, 
        N494, I196_un1_Y, \next_off_div[19] , N498, N499, 
        \nsum_adj_11[17] , I_49_0, \sum_adj[12]_net_1 , N643, 
        I204_un1_Y, N595, N530, \next_off_div[22] , \next_off_div[4] , 
        \nsum_adj_11[20] , I_59_0, \nsum_adj_11[19] , I_56_0, N_2, 
        \DWACT_FINC_E[29] , \DWACT_FINC_E[13] , \DWACT_FINC_E[33] , 
        \DWACT_FINC_E[34] , \DWACT_FINC_E[2] , \DWACT_FINC_E[5] , 
        \DWACT_FINC_E[15] , N_3, \DWACT_FINC_E[28] , 
        \DWACT_FINC_E[16] , N_4, N_5, \DWACT_FINC_E[14] , N_6, 
        \DWACT_FINC_E[9] , \DWACT_FINC_E[12] , N_7, \DWACT_FINC_E[10] , 
        \DWACT_FINC_E[0] , N_8, \DWACT_FINC_E[11] , N_9, N_10, N_11, 
        \DWACT_FINC_E[8] , N_12, N_14, N_15, \DWACT_FINC_E[3] , N_17, 
        GND, VCC;
    
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I59_Y (.A(sum_1_0), .B(
        off_div[17]), .C(N432), .Y(N505));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_2 (.A(N482), .B(
        ADD_32x32_fast_I258_Y_0), .C(N551), .Y(ADD_32x32_fast_I258_Y_2)
        );
    NOR2 \off_div_RNI02RJ[30]  (.A(off_div[30]), .B(off_div[29]), .Y(
        next_off_div_2_sqmuxa_5));
    DFN1C0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[0]_net_1 ));
    DFN1E0C0 \off_div[29]  (.D(\next_off_div[29] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[29]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y_0 (.A(N555), .B(N563), 
        .Y(ADD_32x32_fast_I264_Y_0));
    DFN1E0C0 \off_div[26]  (.D(\next_off_div[26] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[26]));
    XOR2 \sum_adj_RNIJMNB[18]  (.A(\sum_adj[18]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[10] ));
    NOR2 \off_div_RNISSPJ[22]  (.A(off_div[22]), .B(off_div[24]), .Y(
        un1_off_divlto31_8));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I247_Y (.A(I247_un1_Y), .B(
        N651), .Y(N796));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I108_Y (.A(N496), .B(N492), 
        .Y(N557));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I47_Y (.A(off_div[23]), .B(
        off_div[22]), .C(sum_0_0), .Y(N493));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I3_P0N (.A(sum_2_0), .B(
        \sum_adj[11]_net_1 ), .C(off_div[3]), .Y(N393));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I165_Y (.A(N489), .B(N493), 
        .C(N562), .Y(N620));
    XNOR2 un13_nsum_adj_I_49 (.A(sum_17), .B(N_8), .Y(I_49_0));
    NOR3 un13_nsum_adj_I_10 (.A(sum_1_d0), .B(sum_0_d0), .C(sum_2_d0), 
        .Y(\DWACT_FINC_E[0] ));
    DFN1E0C0 \off_div[31]  (.D(\next_off_div[31] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[31]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I149_Y (.A(N537), .B(N533), 
        .Y(N598));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I135_Y (.A(N519), .B(N523), 
        .Y(N584));
    AND3 un13_nsum_adj_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[6] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I147_Y (.A(N535), .B(N531), 
        .Y(N596));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I121_Y (.A(N505), .B(N509), 
        .Y(N570));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I272_Y_0 (.A(
        ADD_32x32_fast_I272_un1_Y_0), .B(N638), .C(N637), .Y(
        ADD_32x32_fast_I272_Y_0));
    NOR3A \off_div_RNIURF71[14]  (.A(un1_off_divlto31_4), .B(
        off_div[14]), .C(off_div[15]), .Y(un1_off_divlto31_13));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I173_Y (.A(N562), .B(N570), 
        .Y(N628));
    MX2 \sum_adj_RNO[9]  (.A(sum_9), .B(I_26_0), .S(sum_1_0), .Y(
        \nsum_adj_11[9] ));
    XA1 \off_div_RNO[22]  (.A(N767), .B(ADD_32x32_fast_I312_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[22] ));
    NOR2 \off_div_RNIPNNJ[13]  (.A(off_div[12]), .B(off_div[13]), .Y(
        un1_off_divlto31_2));
    XOR2 \sum_adj_RNIDHOB[21]  (.A(\sum_adj[21]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[13] ));
    DFN1E1C0 \sum_adj[23]  (.D(\nsum_adj_11[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[23]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I203_Y (.A(N594), .B(N601), 
        .C(N593), .Y(N659));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I155_Y (.A(N483), .B(
        ADD_32x32_fast_I155_Y_0), .C(N552), .Y(N610));
    NOR2 un13_nsum_adj_I_57 (.A(sum_19), .B(sum_18), .Y(
        \DWACT_FINC_E[14] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I86_Y (.A(N389), .B(N393), .C(
        N392), .Y(N532));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I200_Y (.A(N597), .B(N590), 
        .C(N589), .Y(N655));
    MX2 \sum_adj_RNO[15]  (.A(sum_15), .B(I_43_0), .S(sum_1_0), .Y(
        \nsum_adj_11[15] ));
    XNOR2 un13_nsum_adj_I_53 (.A(sum_18), .B(N_7), .Y(I_53_0));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I315_Y_0 (.A(off_div[25]), 
        .B(sum_39), .Y(ADD_32x32_fast_I315_Y_0));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I84_Y (.A(N392), .B(
        off_div[4]), .C(\un1_sum_adj[4] ), .Y(N530));
    NOR3B un13_nsum_adj_I_45 (.A(\DWACT_FINC_E[10] ), .B(
        \DWACT_FINC_E[6] ), .C(sum_15), .Y(N_9));
    OR2 \off_div_RNIUMME8[31]  (.A(un1_off_div), .B(off_div[31]), .Y(
        next_off_div37));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I130_Y (.A(N518), .B(N515), 
        .C(N514), .Y(N579));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I266_Y (.A(
        ADD_32x32_fast_I266_un1_Y_0), .B(N657), .C(
        ADD_32x32_fast_I266_Y_0), .Y(N765));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I118_Y (.A(N506), .B(N503), 
        .C(N502), .Y(N567));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I273_un1_Y_0 (.A(N590), .B(
        N598), .C(\un1_sum_adj[0] ), .Y(ADD_32x32_fast_I273_un1_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I69_Y (.A(off_div[12]), .B(
        \un1_sum_adj[12] ), .C(N417), .Y(N515));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I262_Y_0 (.A(N551), .B(N559), 
        .Y(ADD_32x32_fast_I262_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I202_Y (.A(N592), .B(N599), 
        .C(N591), .Y(N657));
    MX2 \sum_adj_RNO[16]  (.A(sum_16), .B(I_46_0), .S(sum_1_0), .Y(
        \nsum_adj_11[16] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I309_Y_0 (.A(off_div[19]), 
        .B(sum_39), .Y(ADD_32x32_fast_I309_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I184_un1_Y (.A(N581), .B(
        N574), .Y(I184_un1_Y));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I5_P0N (.A(\un1_sum_adj[5] ), 
        .B(off_div[5]), .Y(N399));
    MX2 \off_div_RNO[3]  (.A(next_off_div_0_sqmuxa), .B(
        \un1_off_div_1[3] ), .S(\state_d_0[2] ), .Y(\next_off_div[3] ));
    AND3 un13_nsum_adj_I_69 (.A(\DWACT_FINC_E[29] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[33] ), .Y(N_2));
    NOR3A \off_div_RNISRH71[18]  (.A(un1_off_divlto31_6), .B(
        off_div[19]), .C(off_div[18]), .Y(un1_off_divlto31_14));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I76_Y (.A(N404), .B(
        off_div[8]), .C(\un1_sum_adj[8] ), .Y(N522));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I4_G0N (.A(\un1_sum_adj[4] )
        , .B(off_div[4]), .Y(N395));
    XOR2 \sum_adj_RNIUU1K[14]  (.A(\sum_adj[14]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[6] ));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I1_P0N (.A(\un1_sum_adj[1] ), 
        .B(off_div[1]), .Y(N387));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I13_G0N (.A(
        \un1_sum_adj[13] ), .B(off_div[13]), .Y(N422));
    DFN1E0C0 \off_div[15]  (.D(\next_off_div[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[15]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I150_Y (.A(I150_un1_Y), .B(
        N534), .Y(N599));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I144_Y (.A(N532), .B(N529), 
        .C(N528), .Y(N593));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I74_Y (.A(N407), .B(N411), .C(
        N410), .Y(N520));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I50_Y (.A(off_div[20]), .B(
        off_div[21]), .C(sum_0_0), .Y(N496));
    DFN1E0C0 \off_div[13]  (.D(\next_off_div[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[13]));
    MX2 \sum_adj_RNO[20]  (.A(sum_20), .B(I_59_0), .S(sum_1_0), .Y(
        \nsum_adj_11[20] ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I293_Y_0 (.A(sum_1_0), .B(
        \sum_adj[11]_net_1 ), .C(off_div[3]), .Y(
        ADD_32x32_fast_I293_Y_0));
    AND2 un13_nsum_adj_I_44 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[9] ), .Y(\DWACT_FINC_E[10] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I272_un1_Y_0 (.A(N538), .B(
        N654), .Y(ADD_32x32_fast_I272_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I265_un1_Y (.A(
        ADD_32x32_fast_I265_un1_Y_0), .B(N802), .Y(I265_un1_Y));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I319_Y_0 (.A(off_div[29]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I319_Y_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I265_Y_0 (.A(N557), .B(N565), 
        .Y(ADD_32x32_fast_I265_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I179_Y (.A(N576), .B(N568), 
        .Y(N634));
    AND3 un13_nsum_adj_I_39 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[8] ), .Y(N_11));
    XA1 \off_div_RNO[24]  (.A(N763), .B(ADD_32x32_fast_I314_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[24] ));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I309_Y (.A(I270_un1_Y), .B(
        ADD_32x32_fast_I270_Y_0), .C(ADD_32x32_fast_I309_Y_0), .Y(
        \un1_off_div_1[19] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I177_Y (.A(N566), .B(N574), 
        .Y(N632));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I51_Y (.A(off_div[20]), .B(
        off_div[21]), .C(sum_0_0), .Y(N497));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I308_Y_0 (.A(off_div[18]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I308_Y_0));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I2_P0N (.A(sum_2_0), .B(
        \sum_adj[10]_net_1 ), .C(off_div[2]), .Y(N390));
    NOR2 \state_RNIRG6H_2[0]  (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(pwm_rdy));
    OA1 \off_div_RNIE0NM[1]  (.A(off_div[0]), .B(off_div[1]), .C(
        off_div[2]), .Y(un5lt4));
    DFN1E0P0 \off_div[7]  (.D(\next_off_div[7] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[7]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I196_Y (.A(I196_un1_Y), .B(
        N585), .Y(N651));
    NOR3 un13_nsum_adj_I_29 (.A(sum_7), .B(sum_6), .C(sum_8), .Y(
        \DWACT_FINC_E[5] ));
    NOR2A \state_RNIRG6H_0[0]  (.A(\state[1]_net_1 ), .B(
        \state[0]_net_1 ), .Y(\state_d_0[2] ));
    XNOR2 un13_nsum_adj_I_65 (.A(sum_22), .B(N_3), .Y(I_65_0));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I268_Y (.A(I230_un1_Y), .B(
        N629), .C(I268_un1_Y), .Y(N769));
    DFN1E0C0 \off_div[9]  (.D(\next_off_div[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[9]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I37_Y (.A(off_div[28]), .B(
        off_div[27]), .C(sum_2_0), .Y(N483));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I186_Y (.A(N583), .B(N576), 
        .C(N575), .Y(N641));
    DFN1E0C0 \off_div[11]  (.D(\next_off_div[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[11]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I145_Y (.A(N533), .B(N529), 
        .Y(N594));
    DFN1E1C0 \sum_adj[18]  (.D(\nsum_adj_11[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[18]_net_1 ));
    MX2 un1_off_div_1_0_0_ADD_32x32_fast_I92_Y (.A(sum_1_0), .B(
        off_div[0]), .S(\sum_adj[8]_net_1 ), .Y(N538));
    XA1 \off_div_RNO[13]  (.A(N787), .B(ADD_32x32_fast_I303_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[13] ));
    MX2 \sum_adj_RNO[21]  (.A(sum_21), .B(I_62_0), .S(sum_1_0), .Y(
        \nsum_adj_11[21] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I318_Y_0 (.A(off_div[28]), 
        .B(sum_39), .Y(ADD_32x32_fast_I318_Y_0));
    XNOR2 un13_nsum_adj_I_35 (.A(sum_12), .B(N_13), .Y(I_35_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I191_Y (.A(N588), .B(N580), 
        .Y(N646));
    MX2 \sum_adj_RNO[22]  (.A(sum_22), .B(I_65_0), .S(sum_1_0), .Y(
        \nsum_adj_11[22] ));
    MX2 \off_div_RNO[15]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[15] ), .S(\state_d_0[2] ), .Y(
        \next_off_div[15] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y (.A(
        ADD_32x32_fast_I258_un1_Y_0), .B(N781), .C(
        ADD_32x32_fast_I258_Y_3), .Y(N749));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I14_P0N (.A(sum_2_0), .B(
        \sum_adj[22]_net_1 ), .C(off_div[14]), .Y(N426));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I122_Y (.A(N510), .B(N507), 
        .C(N506), .Y(N571));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I89_Y (.A(N387), .B(N390), 
        .Y(N535));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I262_Y_1 (.A(N618), .B(N633), 
        .C(ADD_32x32_fast_I262_Y_0), .Y(ADD_32x32_fast_I262_Y_1));
    AND3 un13_nsum_adj_I_64 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[16] ), .Y(N_3));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I265_Y (.A(I224_un1_Y), .B(
        ADD_32x32_fast_I265_Y_0), .C(I265_un1_Y), .Y(N763));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I181_Y (.A(N578), .B(N570), 
        .Y(N636));
    NOR2A un13_nsum_adj_I_25 (.A(\DWACT_FINC_E[4] ), .B(sum_8), .Y(
        N_16));
    DFN1E1C0 \sum_adj[9]  (.D(\nsum_adj_11[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[9]_net_1 ));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I60_Y (.A(N428), .B(sum_1_0), 
        .C(off_div[16]), .Y(N506));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I307_Y (.A(I238_un1_Y), .B(
        ADD_32x32_fast_I272_Y_0), .C(ADD_32x32_fast_I307_Y_0), .Y(
        \un1_off_div_1[17] ));
    AND3 un13_nsum_adj_I_51 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[28] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I174_Y (.A(N571), .B(N564), 
        .C(N563), .Y(N629));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I140_Y (.A(N528), .B(N525), 
        .C(N524), .Y(N589));
    DFN1E1C0 \sum_adj[11]  (.D(\nsum_adj_11[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[11]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y_1 (.A(N620), .B(N635), 
        .C(ADD_32x32_fast_I263_Y_0), .Y(ADD_32x32_fast_I263_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I246_Y (.A(N650), .B(N599), 
        .C(N649), .Y(N793));
    XA1 \off_div_RNO[27]  (.A(N757), .B(ADD_32x32_fast_I317_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[27] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I291_Y_0 (.A(off_div[1]), .B(
        \un1_sum_adj[1] ), .Y(ADD_32x32_fast_I291_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I249_un1_Y (.A(N590), .B(
        N598), .C(\un1_sum_adj[0] ), .Y(I249_un1_Y));
    NOR2B \off_div_RNIUTOJ[19]  (.A(off_div[19]), .B(off_div[20]), .Y(
        un5lto20_1));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I13_P0N (.A(\un1_sum_adj[13] )
        , .B(off_div[13]), .Y(N423));
    AND3 un13_nsum_adj_I_48 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[11] ), .Y(N_8));
    DFN1E0C0 \off_div[25]  (.D(\next_off_div[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[25]));
    XA1 \off_div_RNO[1]  (.A(N538), .B(ADD_32x32_fast_I291_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[1] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I61_Y (.A(N432), .B(N429), 
        .Y(N507));
    NOR2B un13_nsum_adj_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_13));
    DFN1E1C0 \sum_adj[22]  (.D(\nsum_adj_11[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[22]_net_1 ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I79_Y (.A(off_div[6]), .B(
        \un1_sum_adj[6] ), .C(N405), .Y(N525));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I150_un1_Y (.A(N535), .B(
        N538), .Y(I150_un1_Y));
    OA1 \off_div_RNIH9KL2[10]  (.A(un5lto9), .B(un5lt9), .C(
        off_div[10]), .Y(un5lt14));
    DFN1E0C0 \off_div[23]  (.D(\next_off_div[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[23]));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I304_Y_0 (.A(sum_0_0), .B(
        \sum_adj[22]_net_1 ), .C(off_div[14]), .Y(
        ADD_32x32_fast_I304_Y_0));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I298_Y_0 (.A(off_div[8]), .B(
        \un1_sum_adj[8] ), .Y(ADD_32x32_fast_I298_Y_0));
    XA1 \off_div_RNO[9]  (.A(N799), .B(ADD_32x32_fast_I299_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[9] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y_1 (.A(N622), .B(N637), 
        .C(ADD_32x32_fast_I264_Y_0), .Y(ADD_32x32_fast_I264_Y_1));
    GND GND_i (.Y(GND));
    AND3 un13_nsum_adj_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E[4] ));
    DFN1E1C0 \sum_adj[14]  (.D(\nsum_adj_11[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[14]_net_1 ));
    OR2 \off_div_RNIPQ4F[3]  (.A(off_div[4]), .B(off_div[3]), .Y(
        un5lto4));
    NOR3B \off_div_RNI30B61[31]  (.A(\state[0]_net_1 ), .B(
        next_off_div_2_sqmuxa_1), .C(off_div[31]), .Y(
        next_off_div_2_sqmuxa_6));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I138_Y (.A(N526), .B(N523), 
        .C(N522), .Y(N587));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y (.A(
        ADD_32x32_fast_I259_un1_Y_0), .B(N784), .C(
        ADD_32x32_fast_I259_Y_3), .Y(N751));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I43_Y (.A(off_div[25]), .B(
        off_div[24]), .C(sum_0_0), .Y(N489));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I123_Y (.A(N511), .B(N507), 
        .Y(N572));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I175_Y (.A(N564), .B(N572), 
        .Y(N630));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I106_Y (.A(N490), .B(N494), 
        .Y(N555));
    MX2 \sum_adj_RNO[10]  (.A(sum_10), .B(I_28_0), .S(sum_1_0), .Y(
        \nsum_adj_11[10] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I11_G0N (.A(
        \un1_sum_adj[11] ), .B(off_div[11]), .Y(N416));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I314_Y_0 (.A(off_div[24]), 
        .B(sum_39), .Y(ADD_32x32_fast_I314_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I271_un1_Y_0 (.A(N586), .B(
        N594), .C(N601), .Y(ADD_32x32_fast_I271_un1_Y_0));
    DFN1E0C0 \off_div[21]  (.D(\next_off_div[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[21]));
    XA1 \off_div_RNO[11]  (.A(N793), .B(ADD_32x32_fast_I301_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[11] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I42_Y (.A(off_div[24]), .B(
        off_div[25]), .C(sum_0_0), .Y(N488));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y (.A(
        ADD_32x32_fast_I263_un1_Y_0), .B(N796), .C(
        ADD_32x32_fast_I263_Y_1), .Y(N759));
    OA1 \off_div_RNI3NCO5[16]  (.A(off_div[16]), .B(un5lt16), .C(
        un5lto20_2), .Y(un5lt31));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I248_Y (.A(N654), .B(N538), 
        .C(N653), .Y(N799));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I301_Y_0 (.A(off_div[11]), 
        .B(\un1_sum_adj[11] ), .Y(ADD_32x32_fast_I301_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y (.A(
        ADD_32x32_fast_I260_un1_Y_0), .B(N787), .C(
        ADD_32x32_fast_I260_Y_2), .Y(N753));
    AND3 un13_nsum_adj_I_68 (.A(\DWACT_FINC_E[34] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[29] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I306_Y_0 (.A(off_div[16]), 
        .B(sum_39), .Y(ADD_32x32_fast_I306_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I155_Y_0 (.A(off_div[29]), .B(
        off_div[30]), .C(sum_0_0), .Y(ADD_32x32_fast_I155_Y_0));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I80_Y (.A(N398), .B(
        off_div[6]), .C(\un1_sum_adj[6] ), .Y(N526));
    DFN1E1C0 \sum_adj[13]  (.D(\nsum_adj_11[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[13]_net_1 ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I265_un1_Y_0 (.A(N624), .B(
        N640), .Y(ADD_32x32_fast_I265_un1_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I262_Y (.A(
        ADD_32x32_fast_I262_un1_Y_0), .B(N793), .C(
        ADD_32x32_fast_I262_Y_1), .Y(N757));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I170_Y (.A(N567), .B(N560), 
        .C(N559), .Y(N625));
    DFN1E0C0 \off_div[5]  (.D(\next_off_div[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[5]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I7_G0N (.A(\un1_sum_adj[7] )
        , .B(off_div[7]), .Y(N404));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I57_Y (.A(off_div[17]), .B(
        off_div[18]), .C(sum_0_0), .Y(N503));
    XOR2 \state_RNO[1]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 ), 
        .Y(N_311_i));
    NOR3 un13_nsum_adj_I_18 (.A(sum_5), .B(sum_4), .C(sum_3), .Y(
        \DWACT_FINC_E[2] ));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I308_Y (.A(I236_un1_Y), .B(
        ADD_32x32_fast_I271_Y_0), .C(ADD_32x32_fast_I308_Y_0), .Y(
        \un1_off_div_1[18] ));
    MX2 \sum_adj_RNO[11]  (.A(sum_11), .B(I_32_0), .S(sum_1_0), .Y(
        \nsum_adj_11[11] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I321_Y_0 (.A(off_div[31]), 
        .B(sum_39), .Y(ADD_32x32_fast_I321_Y_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I116_Y (.A(N504), .B(N500), 
        .Y(N565));
    NOR2 un13_nsum_adj_I_38 (.A(sum_12), .B(sum_13), .Y(
        \DWACT_FINC_E[8] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I311_Y_0 (.A(off_div[21]), 
        .B(sum_39), .Y(ADD_32x32_fast_I311_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I269_Y_0 (.A(N647), .B(N632), 
        .C(N631), .Y(ADD_32x32_fast_I269_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I81_Y (.A(off_div[6]), .B(
        \un1_sum_adj[6] ), .C(N399), .Y(N527));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I245_Y (.A(N648), .B(N663), 
        .C(N647), .Y(N790));
    MX2 \sum_adj_RNO[12]  (.A(sum_12), .B(I_35_0), .S(sum_1_0), .Y(
        \nsum_adj_11[12] ));
    NOR2B \off_div_RNIUVJ71[23]  (.A(next_off_div_2_sqmuxa_2), .B(
        un1_off_divlto31_9), .Y(next_off_div_2_sqmuxa_7));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I316_Y_0 (.A(off_div[26]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I316_Y_0));
    XNOR2 un13_nsum_adj_I_46 (.A(sum_16), .B(N_9), .Y(I_46_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I70_Y (.A(N413), .B(N417), .C(
        N416), .Y(N516));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I192_Y (.A(N589), .B(N582), 
        .C(N581), .Y(N647));
    XNOR2 un13_nsum_adj_I_28 (.A(sum_10), .B(N_15), .Y(I_28_0));
    DFN1E0C0 \off_div[30]  (.D(\next_off_div[30] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[30]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I129_Y (.A(N513), .B(N517), 
        .Y(N578));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I182_Y (.A(N579), .B(N572), 
        .C(N571), .Y(N637));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I127_Y (.A(N511), .B(N515), 
        .Y(N576));
    XOR2 \sum_adj_RNIKNNB[19]  (.A(\sum_adj[19]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[11] ));
    VCC VCC_i (.Y(VCC));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I249_Y (.A(I249_un1_Y), .B(
        N655), .Y(N802));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I0_G0N (.A(off_div[0]), .B(
        sum_39), .Y(N383));
    NOR3C \off_div_RNITFNM[5]  (.A(off_div[5]), .B(off_div[7]), .C(
        off_div[6]), .Y(un5lto7_1));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I196_un1_Y (.A(N593), .B(
        N586), .Y(I196_un1_Y));
    AO1C \state_RNI5VA5I_0[1]  (.A(un5lt31), .B(
        next_off_div_2_sqmuxa_11), .C(\state[1]_net_1 ), .Y(
        un1_state_2));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I45_Y (.A(off_div[24]), .B(
        off_div[23]), .C(sum_0_0), .Y(N491));
    AND3 un13_nsum_adj_I_52 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[12] ), .Y(N_7));
    NOR3A \off_div_RNIEBF71[11]  (.A(un1_off_divlto31_2), .B(
        off_div[11]), .C(off_div[10]), .Y(un1_off_divlto31_12));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I111_Y (.A(N495), .B(N499), 
        .Y(N560));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I71_Y (.A(off_div[10]), .B(
        \un1_sum_adj[10] ), .C(N417), .Y(N517));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I9_G0N (.A(\un1_sum_adj[9] )
        , .B(off_div[9]), .Y(N410));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I228_un1_Y (.A(N643), .B(
        N628), .Y(I228_un1_Y));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I307_Y_0 (.A(off_div[17]), 
        .B(sum_39), .Y(ADD_32x32_fast_I307_Y_0));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I2_G0N (.A(sum_1_0), .B(
        \sum_adj[10]_net_1 ), .C(off_div[2]), .Y(N389));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I148_Y (.A(N536), .B(N533), 
        .C(N532), .Y(N597));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I48_Y (.A(off_div[21]), .B(
        off_div[22]), .C(sum_0_0), .Y(N494));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I260_un1_Y_0 (.A(N614), .B(
        N630), .Y(ADD_32x32_fast_I260_un1_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I268_un1_Y (.A(N630), .B(
        N646), .C(N661), .Y(I268_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_3 (.A(N612), .B(N627), 
        .C(ADD_32x32_fast_I259_Y_2), .Y(ADD_32x32_fast_I259_Y_3));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I266_un1_Y_0 (.A(N642), .B(
        N626), .Y(ADD_32x32_fast_I266_un1_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I67_Y (.A(off_div[12]), .B(
        \un1_sum_adj[12] ), .C(N423), .Y(N513));
    XNOR2 un13_nsum_adj_I_70 (.A(sum_23), .B(N_2), .Y(I_70_0));
    NOR3A un13_nsum_adj_I_66 (.A(\DWACT_FINC_E[15] ), .B(sum_21), .C(
        sum_22), .Y(\DWACT_FINC_E[33] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I193_Y (.A(N582), .B(N590), 
        .Y(N648));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I5_G0N (.A(\un1_sum_adj[5] )
        , .B(off_div[5]), .Y(N398));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I317_Y_0 (.A(off_div[27]), 
        .B(sum_39), .Y(ADD_32x32_fast_I317_Y_0));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y_1 (.A(N486), .B(N482), 
        .C(N555), .Y(ADD_32x32_fast_I260_Y_1));
    XOR2 \sum_adj_RNIVV1K[15]  (.A(\sum_adj[15]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[7] ));
    NOR2 \off_div_RNI12QJ[25]  (.A(off_div[26]), .B(off_div[25]), .Y(
        un1_off_divlto31_9));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I243_Y (.A(N644), .B(N659), 
        .C(N643), .Y(N784));
    NOR2 \off_div_RNINNPJ[20]  (.A(off_div[20]), .B(off_div[21]), .Y(
        un1_off_divlto31_6));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I296_Y_0 (.A(off_div[6]), .B(
        \un1_sum_adj[6] ), .Y(ADD_32x32_fast_I296_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I183_Y (.A(N572), .B(N580), 
        .Y(N638));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I157_Y_1 (.A(
        ADD_32x32_fast_I157_Y_0), .B(N485), .Y(ADD_32x32_fast_I157_Y_1)
        );
    MX2 \sum_adj_RNO[8]  (.A(sum_8), .B(I_23_2), .S(sum_1_0), .Y(
        \nsum_adj_11[8] ));
    XA1 \off_div_RNO[6]  (.A(N659), .B(ADD_32x32_fast_I296_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[6] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I124_Y (.A(N512), .B(N509), 
        .C(N508), .Y(N573));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I273_Y_0 (.A(
        ADD_32x32_fast_I273_un1_Y_0), .B(N640), .C(N639), .Y(
        ADD_32x32_fast_I273_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I157_Y_0 (.A(off_div[28]), .B(
        off_div[29]), .C(sum_2_0), .Y(ADD_32x32_fast_I157_Y_0));
    NOR2 \off_div_RNITTPJ[23]  (.A(off_div[23]), .B(off_div[24]), .Y(
        next_off_div_2_sqmuxa_2));
    NOR3B un13_nsum_adj_I_36 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .C(sum_12), .Y(N_12));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I242_Y (.A(N642), .B(N657), 
        .C(N641), .Y(N781));
    XOR2 \sum_adj_RNI218E[8]  (.A(\sum_adj[8]_net_1 ), .B(sum_2_0), .Y(
        \un1_sum_adj[0] ));
    DFN1E0C0 \off_div[1]  (.D(\next_off_div[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[1]));
    NOR2 un13_nsum_adj_I_47 (.A(sum_15), .B(sum_16), .Y(
        \DWACT_FINC_E[11] ));
    XA1 \off_div_RNO[8]  (.A(N802), .B(ADD_32x32_fast_I298_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[8] ));
    NOR2B \off_div_RNI58L71[30]  (.A(un1_off_divlto31_10), .B(
        next_off_div_2_sqmuxa_5), .Y(next_off_div_2_sqmuxa_8));
    XNOR2 un13_nsum_adj_I_26 (.A(sum_9), .B(N_16), .Y(I_26_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I102_Y (.A(N490), .B(N486), 
        .Y(N551));
    XNOR2 un13_nsum_adj_I_43 (.A(sum_15), .B(N_10), .Y(I_43_0));
    MX2 \off_div_RNO[19]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[19] ), .S(\state_d_0[2] ), .Y(
        \next_off_div[19] ));
    DFN1E0C0 \off_div[10]  (.D(\next_off_div[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[10]));
    MX2 \off_div_RNO[10]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[10] ), .S(\state_d_0[2] ), .Y(
        \next_off_div[10] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I125_Y (.A(N513), .B(N509), 
        .Y(N574));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y_0 (.A(N553), .B(N561), 
        .Y(ADD_32x32_fast_I263_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I178_Y (.A(N575), .B(N568), 
        .C(N567), .Y(N633));
    DFN1E1C0 \sum_adj[12]  (.D(\nsum_adj_11[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[12]_net_1 ));
    NOR3 un13_nsum_adj_I_50 (.A(sum_16), .B(sum_15), .C(sum_17), .Y(
        \DWACT_FINC_E[12] ));
    MX2 \sum_adj_RNO[17]  (.A(sum_17), .B(I_49_0), .S(sum_1_0), .Y(
        \nsum_adj_11[17] ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I297_Y (.A(\un1_sum_adj[7] ), 
        .B(off_div[7]), .C(N657), .Y(\un1_off_div_1[7] ));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I269_un1_Y (.A(N632), .B(
        N648), .C(N663), .Y(I269_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I136_Y (.A(N524), .B(N521), 
        .C(N520), .Y(N585));
    XA1 \off_div_RNO[16]  (.A(N779), .B(ADD_32x32_fast_I306_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[16] ));
    XOR2 \sum_adj_RNITT1K[13]  (.A(\sum_adj[13]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[5] ));
    NOR3A \off_div_RNIMA781[29]  (.A(un1_off_divlto31_0), .B(
        off_div[29]), .C(un5lto9), .Y(un1_off_divlto31_17));
    MX2 \off_div_RNO[0]  (.A(next_off_div_0_sqmuxa), .B(
        \un1_off_div_1[0] ), .S(\state_d_0[2] ), .Y(\next_off_div[0] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I199_Y (.A(N596), .B(N588), 
        .Y(N654));
    XA1 \off_div_RNO[23]  (.A(N765), .B(ADD_32x32_fast_I313_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[23] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I264_un1_Y_0 (.A(N622), .B(
        N638), .Y(ADD_32x32_fast_I264_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I87_Y (.A(N390), .B(N393), 
        .Y(N533));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I189_Y (.A(N578), .B(N586), 
        .Y(N644));
    XOR2 \sum_adj_RNISS1K[12]  (.A(\sum_adj[12]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[4] ));
    MX2 \off_div_RNO[18]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[18] ), .S(\state_d_0[2] ), .Y(
        \next_off_div[18] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I38_Y (.A(off_div[27]), .B(
        off_div[26]), .C(sum_2_0), .Y(N484));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I187_Y (.A(N576), .B(N584), 
        .Y(N642));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I273_Y (.A(N655), .B(N640), 
        .C(ADD_32x32_fast_I273_Y_0), .Y(N779));
    NOR3 un13_nsum_adj_I_67 (.A(sum_1_d0), .B(sum_0_d0), .C(sum_2_d0), 
        .Y(\DWACT_FINC_E[34] ));
    XA1 \off_div_RNO[25]  (.A(N761), .B(ADD_32x32_fast_I315_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[25] ));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I112_Y (.A(N496), .B(N500), 
        .Y(N561));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I14_G0N (.A(sum_2_0), .B(
        \sum_adj[22]_net_1 ), .C(off_div[14]), .Y(N425));
    DFN1E0C0 \off_div[12]  (.D(\next_off_div[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[12]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I271_Y_0 (.A(
        ADD_32x32_fast_I271_un1_Y_0), .B(N636), .C(N635), .Y(
        ADD_32x32_fast_I271_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I161_Y (.A(
        ADD_32x32_fast_I161_Y_0), .B(N558), .Y(N616));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I103_Y (.A(N491), .B(N487), 
        .Y(N552));
    DFN1E0C0 \off_div[0]  (.D(\next_off_div[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[0]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I131_Y (.A(N515), .B(N519), 
        .Y(N580));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I120_Y (.A(N508), .B(N505), 
        .C(N504), .Y(N569));
    NOR2A un13_nsum_adj_I_63 (.A(\DWACT_FINC_E[15] ), .B(sum_21), .Y(
        \DWACT_FINC_E[16] ));
    NOR2 \off_div_RNI10OJ[16]  (.A(off_div[17]), .B(off_div[16]), .Y(
        un1_off_divlto31_4));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I46_Y (.A(off_div[22]), .B(
        off_div[23]), .C(sum_0_0), .Y(N492));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I300_Y_0 (.A(off_div[10]), 
        .B(\un1_sum_adj[10] ), .Y(ADD_32x32_fast_I300_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I77_Y (.A(off_div[8]), .B(
        \un1_sum_adj[8] ), .C(N405), .Y(N523));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I44_Y (.A(off_div[23]), .B(
        off_div[24]), .C(sum_0_0), .Y(N490));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y_2 (.A(N614), .B(N629), 
        .C(ADD_32x32_fast_I260_Y_1), .Y(ADD_32x32_fast_I260_Y_2));
    DFN1E1C0 \sum_adj[20]  (.D(\nsum_adj_11[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[20]_net_1 ));
    OR3 \off_div_RNIIFF71[11]  (.A(off_div[12]), .B(off_div[11]), .C(
        un5lto14_1), .Y(un5lto14_2));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I53_Y (.A(off_div[19]), .B(
        off_div[20]), .C(sum_0_0), .Y(N499));
    MX2 \off_div_RNO[5]  (.A(next_off_div_0_sqmuxa), .B(
        \un1_off_div_1[5] ), .S(\state_d_0[2] ), .Y(\next_off_div[5] ));
    XNOR2 un13_nsum_adj_I_37 (.A(sum_13), .B(N_12), .Y(I_37_0));
    XA1 \off_div_RNO[2]  (.A(N601), .B(ADD_32x32_fast_I292_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[2] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I6_G0N (.A(\un1_sum_adj[6] )
        , .B(off_div[6]), .Y(N401));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I247_un1_Y (.A(N586), .B(
        N594), .C(N601), .Y(I247_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I151_Y (.A(N537), .B(
        \un1_sum_adj[0] ), .C(N536), .Y(N601));
    DFN1E0C0 \off_div[6]  (.D(\next_off_div[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[6]));
    NOR3 un13_nsum_adj_I_33 (.A(sum_10), .B(sum_9), .C(sum_11), .Y(
        \DWACT_FINC_E[7] ));
    DFN1E1C0 \sum_adj[17]  (.D(\nsum_adj_11[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[17]_net_1 ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I320_Y_0 (.A(off_div[30]), 
        .B(sum_39), .Y(ADD_32x32_fast_I320_Y_0));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I305_Y (.A(\un1_sum_adj[15] )
        , .B(off_div[15]), .C(N781), .Y(\un1_off_div_1[15] ));
    NOR3A un13_nsum_adj_I_27 (.A(\DWACT_FINC_E[4] ), .B(sum_8), .C(
        sum_9), .Y(N_15));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I310_Y_0 (.A(off_div[20]), 
        .B(sum_39), .Y(ADD_32x32_fast_I310_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I270_Y_0 (.A(N649), .B(N634), 
        .C(N633), .Y(ADD_32x32_fast_I270_Y_0));
    XOR2 \sum_adj_RNI328E[9]  (.A(\sum_adj[9]_net_1 ), .B(sum_2_0), .Y(
        \un1_sum_adj[1] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I230_un1_Y (.A(N645), .B(
        N630), .Y(I230_un1_Y));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I52_Y (.A(off_div[20]), .B(
        off_div[19]), .C(sum_0_0), .Y(N498));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I204_Y (.A(I204_un1_Y), .B(
        N595), .Y(N661));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I263_un1_Y_0 (.A(N620), .B(
        N636), .Y(ADD_32x32_fast_I263_un1_Y_0));
    XOR2 \sum_adj_RNI122K[17]  (.A(\sum_adj[17]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[9] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I194_Y (.A(N591), .B(N584), 
        .C(N583), .Y(N649));
    XNOR2 un13_nsum_adj_I_23 (.A(sum_8), .B(N_17), .Y(I_23_2));
    XNOR2 un13_nsum_adj_I_59 (.A(sum_20), .B(N_5), .Y(I_59_0));
    DFN1E0C0 \off_div[20]  (.D(\next_off_div[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[20]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I113_Y (.A(N497), .B(N501), 
        .Y(N562));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I184_Y (.A(I184_un1_Y), .B(
        N573), .Y(N639));
    NOR3 un13_nsum_adj_I_41 (.A(sum_13), .B(sum_12), .C(sum_14), .Y(
        \DWACT_FINC_E[9] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_0 (.A(off_div[29]), .B(
        off_div[28]), .C(sum_1_0), .Y(ADD_32x32_fast_I259_Y_0));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I294_Y_0 (.A(off_div[4]), .B(
        \un1_sum_adj[4] ), .Y(ADD_32x32_fast_I294_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I236_un1_Y (.A(N651), .B(
        N636), .Y(I236_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I10_G0N (.A(
        \un1_sum_adj[10] ), .B(off_div[10]), .Y(N413));
    XA1 \off_div_RNO[21]  (.A(N769), .B(ADD_32x32_fast_I311_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[21] ));
    DFN1E0C0 \off_div[18]  (.D(\next_off_div[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[18]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I262_un1_Y_0 (.A(N618), .B(
        N634), .Y(ADD_32x32_fast_I262_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I109_Y (.A(N497), .B(N493), 
        .Y(N558));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I146_Y (.A(N534), .B(N531), 
        .C(N530), .Y(N595));
    NOR3C \off_div_RNI10H71[17]  (.A(off_div[18]), .B(off_div[17]), .C(
        un5lto20_1), .Y(un5lto20_2));
    NOR3C \state_RNIP7TV8[0]  (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .C(next_off_div37), .Y(
        next_off_div_0_sqmuxa));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I195_Y (.A(N592), .B(N584), 
        .Y(N650));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I63_Y (.A(N426), .B(N429), 
        .Y(N509));
    NOR3C \off_div_RNITHBU1[5]  (.A(un1_off_divlto31_10), .B(
        un1_off_divlto31_9), .C(un1_off_divlt31), .Y(
        un1_off_divlto31_20));
    NOR3B un13_nsum_adj_I_55 (.A(\DWACT_FINC_E[13] ), .B(
        \DWACT_FINC_E[28] ), .C(sum_18), .Y(N_6));
    DFN1E0C0 \off_div[22]  (.D(\next_off_div[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[22]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I185_Y (.A(N574), .B(N582), 
        .Y(N640));
    NOR2A \state_RNIRG6H_1[0]  (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(state_176_d));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I90_Y (.A(N383), .B(N387), .C(
        N386), .Y(N536));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I55_Y (.A(off_div[18]), .B(
        off_div[19]), .C(sum_0_0), .Y(N501));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I49_Y (.A(off_div[22]), .B(
        off_div[21]), .C(sum_0_0), .Y(N495));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_2 (.A(N484), .B(
        ADD_32x32_fast_I259_Y_0), .C(N553), .Y(ADD_32x32_fast_I259_Y_2)
        );
    XA1 \off_div_RNO[12]  (.A(N790), .B(ADD_32x32_fast_I302_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[12] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I62_Y (.A(N425), .B(N429), .C(
        N428), .Y(N508));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y (.A(
        ADD_32x32_fast_I261_un1_Y_0), .B(N790), .C(
        ADD_32x32_fast_I261_Y_2), .Y(N755));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I141_Y (.A(N529), .B(N525), 
        .Y(N590));
    AND3 un13_nsum_adj_I_61 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[15] ), .Y(N_4));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I36_Y (.A(off_div[27]), .B(
        off_div[28]), .C(sum_2_0), .Y(N482));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I7_P0N (.A(\un1_sum_adj[7] ), 
        .B(off_div[7]), .Y(N405));
    NOR2 \off_div_RNI56QJ[27]  (.A(off_div[27]), .B(off_div[28]), .Y(
        un1_off_divlto31_10));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I58_Y (.A(off_div[17]), .B(
        off_div[16]), .C(sum_0_0), .Y(N504));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I292_Y_0 (.A(sum_0_0), .B(
        \sum_adj[10]_net_1 ), .C(off_div[2]), .Y(
        ADD_32x32_fast_I292_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I91_Y (.A(sum_1_0), .B(
        off_div[0]), .C(N387), .Y(N537));
    DFN1E0C0 \off_div[17]  (.D(\next_off_div[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[17]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I119_Y (.A(N503), .B(N507), 
        .Y(N568));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I190_Y (.A(N587), .B(N580), 
        .C(N579), .Y(N645));
    AND3 un13_nsum_adj_I_54 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[9] ), .C(\DWACT_FINC_E[12] ), .Y(
        \DWACT_FINC_E[13] ));
    MX2 \sum_adj_RNO[23]  (.A(sum_23), .B(I_70_0), .S(sum_1_0), .Y(
        \nsum_adj_11[23] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I117_Y (.A(N505), .B(N501), 
        .Y(N566));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I132_Y (.A(N520), .B(N517), 
        .C(N516), .Y(N581));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I180_Y (.A(N577), .B(N570), 
        .C(N569), .Y(N635));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I128_Y (.A(N516), .B(N513), 
        .C(N512), .Y(N577));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I104_Y (.A(N492), .B(N488), 
        .Y(N553));
    NOR3A un13_nsum_adj_I_31 (.A(\DWACT_FINC_E[6] ), .B(sum_9), .C(
        sum_10), .Y(N_14));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I9_P0N (.A(\un1_sum_adj[9] ), 
        .B(off_div[9]), .Y(N411));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I15_G0N (.A(
        \un1_sum_adj[15] ), .B(off_div[15]), .Y(N428));
    OR2 \off_div_RNIRPNJ[13]  (.A(off_div[13]), .B(off_div[14]), .Y(
        un5lto14_1));
    NOR2 un13_nsum_adj_I_21 (.A(sum_6), .B(sum_7), .Y(
        \DWACT_FINC_E[3] ));
    OR2B \off_div_RNIN9NM[5]  (.A(un5lto4), .B(off_div[5]), .Y(
        un1_off_divlt31));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I295_Y_0 (.A(off_div[5]), .B(
        \un1_sum_adj[5] ), .Y(ADD_32x32_fast_I295_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I159_Y_0 (.A(N483), .B(N487)
        , .Y(ADD_32x32_fast_I159_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I176_Y (.A(N573), .B(N566), 
        .C(N565), .Y(N631));
    NOR2 \off_div_RNIPPPJ[21]  (.A(off_div[21]), .B(off_div[22]), .Y(
        next_off_div_2_sqmuxa_1));
    DFN1E0C0 \off_div[28]  (.D(\next_off_div[28] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[28]));
    NOR2B \off_div_RNIHOO48[11]  (.A(un1_off_divlto31_22), .B(
        un1_off_divlto31_21), .Y(un1_off_div));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I83_Y (.A(off_div[4]), .B(
        \un1_sum_adj[4] ), .C(N399), .Y(N529));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I65_Y (.A(N426), .B(N423), 
        .Y(N511));
    DFN1C0 \state[1]  (.D(N_311_i), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \state[1]_net_1 ));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I15_P0N (.A(\un1_sum_adj[15] )
        , .B(off_div[15]), .Y(N429));
    XA1 \off_div_RNO[31]  (.A(N749), .B(ADD_32x32_fast_I321_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[31] ));
    XA1 \off_div_RNO[14]  (.A(N784), .B(ADD_32x32_fast_I304_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[14] ));
    AND3 un13_nsum_adj_I_42 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[9] ), .Y(N_10));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I163_Y (.A(N560), .B(N552), 
        .Y(N618));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I133_Y (.A(N517), .B(N521), 
        .Y(N582));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I68_Y (.A(N416), .B(
        off_div[12]), .C(\un1_sum_adj[12] ), .Y(N514));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I161_Y_0 (.A(N485), .B(N489)
        , .Y(ADD_32x32_fast_I161_Y_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I114_Y (.A(N502), .B(N498), 
        .Y(N563));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I261_un1_Y_0 (.A(N616), .B(
        N632), .Y(ADD_32x32_fast_I261_un1_Y_0));
    NOR3C \off_div_RNI68KL3[31]  (.A(next_off_div_2_sqmuxa_7), .B(
        next_off_div_2_sqmuxa_6), .C(next_off_div_2_sqmuxa_8), .Y(
        next_off_div_2_sqmuxa_10));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I82_Y (.A(N395), .B(N399), .C(
        N398), .Y(N528));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I171_Y (.A(N560), .B(N568), 
        .Y(N626));
    MX2 \sum_adj_RNO[14]  (.A(sum_14), .B(I_40_0), .S(sum_1_0), .Y(
        \nsum_adj_11[14] ));
    NOR2 \off_div_RNIV05F[7]  (.A(off_div[7]), .B(off_div[6]), .Y(
        un1_off_divlto31_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I40_Y (.A(off_div[25]), .B(
        off_div[26]), .C(sum_0_0), .Y(N486));
    DFN1E1C0 \sum_adj[8]  (.D(\nsum_adj_11[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[8]_net_1 ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I204_un1_Y (.A(N596), .B(
        N538), .Y(I204_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I12_G0N (.A(
        \un1_sum_adj[12] ), .B(off_div[12]), .Y(N419));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I11_P0N (.A(\un1_sum_adj[11] )
        , .B(off_div[11]), .Y(N417));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I73_Y (.A(off_div[10]), .B(
        \un1_sum_adj[10] ), .C(N411), .Y(N519));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I266_Y_0 (.A(N641), .B(N626), 
        .C(N625), .Y(ADD_32x32_fast_I266_Y_0));
    NOR2A \state_RNIRG6H[0]  (.A(\state[1]_net_1 ), .B(
        \state[0]_net_1 ), .Y(\state_d[2] ));
    OR2 \off_div_RNI355F[9]  (.A(off_div[9]), .B(off_div[8]), .Y(
        un5lto9));
    AND3 un13_nsum_adj_I_58 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[14] ), .Y(N_5));
    OA1B \state_RNO[0]  (.A(pwm_enable), .B(\state[1]_net_1 ), .C(
        \state[0]_net_1 ), .Y(\state_ns[0] ));
    DFN1E0C0 \off_div[2]  (.D(\next_off_div[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[2]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I39_Y (.A(off_div[27]), .B(
        off_div[26]), .C(sum_2_0), .Y(N485));
    DFN1E0C0 \off_div[27]  (.D(\next_off_div[27] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[27]));
    MX2 \sum_adj_RNO[18]  (.A(sum_18), .B(I_53_0), .S(sum_1_0), .Y(
        \nsum_adj_11[18] ));
    XOR2 \sum_adj_RNI012K[16]  (.A(\sum_adj[16]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[8] ));
    DFN1E1C0 \sum_adj[15]  (.D(\nsum_adj_11[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[15]_net_1 ));
    NOR2A \off_div_RNI4VA4C[31]  (.A(next_off_div_2_sqmuxa_10), .B(
        next_off_div37), .Y(next_off_div_2_sqmuxa_11));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I41_Y (.A(off_div[26]), .B(
        off_div[25]), .C(sum_0_0), .Y(N487));
    OA1 \off_div_RNIINV64[15]  (.A(un5lt14), .B(un5lto14_2), .C(
        off_div[15]), .Y(un5lt16));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y (.A(
        ADD_32x32_fast_I264_un1_Y_0), .B(N799), .C(
        ADD_32x32_fast_I264_Y_1), .Y(N761));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I72_Y (.A(N410), .B(
        off_div[10]), .C(\un1_sum_adj[10] ), .Y(N518));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I295_Y (.A(
        ADD_32x32_fast_I295_Y_0), .B(N661), .Y(\un1_off_div_1[5] ));
    XA1 \off_div_RNO[29]  (.A(N753), .B(ADD_32x32_fast_I319_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[29] ));
    NOR3C \off_div_RNI2I6N3[11]  (.A(un1_off_divlto31_13), .B(
        un1_off_divlto31_12), .C(un1_off_divlto31_17), .Y(
        un1_off_divlto31_21));
    DFN1E0C0 \off_div[14]  (.D(\next_off_div[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[14]));
    DFN1E1C0 \sum_adj[10]  (.D(\nsum_adj_11[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[10]_net_1 ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I302_Y_0 (.A(off_div[12]), 
        .B(\un1_sum_adj[12] ), .Y(ADD_32x32_fast_I302_Y_0));
    MX2 \off_div_RNO[20]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[20] ), .S(\state_d_0[2] ), .Y(
        \next_off_div[20] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I300_Y (.A(
        ADD_32x32_fast_I300_Y_0), .B(N796), .Y(\un1_off_div_1[10] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I115_Y (.A(N499), .B(N503), 
        .Y(N564));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I258_un1_Y_0 (.A(N610), .B(
        N626), .Y(ADD_32x32_fast_I258_un1_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I142_Y (.A(N530), .B(N527), 
        .C(N526), .Y(N591));
    XNOR2 un13_nsum_adj_I_62 (.A(sum_21), .B(N_4), .Y(I_62_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I56_Y (.A(off_div[18]), .B(
        off_div[17]), .C(sum_0_0), .Y(N502));
    XA1 \off_div_RNO[26]  (.A(N759), .B(ADD_32x32_fast_I316_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[26] ));
    MX2 \sum_adj_RNO[13]  (.A(sum_13), .B(I_37_0), .S(sum_1_0), .Y(
        \nsum_adj_11[13] ));
    DFN1E1C0 \sum_adj[19]  (.D(\nsum_adj_11[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[19]_net_1 ));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I267_un1_Y (.A(N628), .B(
        N644), .C(N659), .Y(I267_un1_Y));
    MX2 \off_div_RNO[17]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[17] ), .S(\state_d_0[2] ), .Y(
        \next_off_div[17] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I54_Y (.A(off_div[19]), .B(
        off_div[18]), .C(sum_0_0), .Y(N500));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I267_Y (.A(I228_un1_Y), .B(
        N627), .C(I267_un1_Y), .Y(N767));
    DFN1E0P0 \off_div[4]  (.D(\next_off_div[4] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[4]));
    XOR2 \sum_adj_RNIFJOB[23]  (.A(\sum_adj[23]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[15] ));
    NOR3B \state_RNIP7TV8_0[0]  (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .C(next_off_div37), .Y(
        next_off_div_1_sqmuxa));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I303_Y_0 (.A(off_div[13]), 
        .B(\un1_sum_adj[13] ), .Y(ADD_32x32_fast_I303_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I169_Y (.A(N566), .B(N558), 
        .Y(N624));
    DFN1E0C0 \off_div[19]  (.D(\next_off_div[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[19]));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I85_Y (.A(off_div[4]), .B(
        \un1_sum_adj[4] ), .C(N393), .Y(N531));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I312_Y_0 (.A(off_div[22]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I312_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I139_Y (.A(N527), .B(N523), 
        .Y(N588));
    XOR2 \sum_adj_RNICGOB[20]  (.A(\sum_adj[20]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[12] ));
    XA1 \off_div_RNO[28]  (.A(N755), .B(ADD_32x32_fast_I318_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[28] ));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I167_Y (.A(N495), .B(N491), 
        .C(N564), .Y(N622));
    DFN1E0C0 \off_div[16]  (.D(\next_off_div[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[16]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I198_Y (.A(N595), .B(N588), 
        .C(N587), .Y(N653));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I137_Y (.A(N521), .B(N525), 
        .Y(N586));
    DFN1E0P0 \off_div[8]  (.D(\next_off_div[8] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[8]));
    XNOR2 un13_nsum_adj_I_32 (.A(sum_11), .B(N_14), .Y(I_32_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I188_Y (.A(N585), .B(N578), 
        .C(N577), .Y(N643));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I16_P0N (.A(off_div[16]), .B(
        sum_2_0), .Y(N432));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I110_Y (.A(N498), .B(N494), 
        .Y(N559));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I88_Y (.A(N386), .B(N390), .C(
        N389), .Y(N534));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0 (.A(off_div[30]), .B(
        off_div[29]), .C(sum_0_0), .Y(ADD_32x32_fast_I258_Y_0));
    AND3 un13_nsum_adj_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_17));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I310_Y (.A(I269_un1_Y), .B(
        ADD_32x32_fast_I269_Y_0), .C(ADD_32x32_fast_I310_Y_0), .Y(
        \un1_off_div_1[20] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y_2 (.A(N616), .B(N631), 
        .C(ADD_32x32_fast_I261_Y_1), .Y(ADD_32x32_fast_I261_Y_2));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I159_Y (.A(N495), .B(N491), 
        .C(ADD_32x32_fast_I159_Y_0), .Y(N614));
    XNOR2 un13_nsum_adj_I_40 (.A(sum_14), .B(N_11), .Y(I_40_0));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I313_Y_0 (.A(off_div[23]), 
        .B(sum_39), .Y(ADD_32x32_fast_I313_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I157_Y (.A(N489), .B(N493), 
        .C(ADD_32x32_fast_I157_Y_1), .Y(N612));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I75_Y (.A(off_div[8]), .B(
        \un1_sum_adj[8] ), .C(N411), .Y(N521));
    NOR3C \off_div_RNIF6ID4[18]  (.A(un1_off_divlto31_15), .B(
        un1_off_divlto31_14), .C(un1_off_divlto31_20), .Y(
        un1_off_divlto31_22));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I293_Y (.A(
        ADD_32x32_fast_I293_Y_0), .B(N599), .Y(\un1_off_div_1[3] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I143_Y (.A(N527), .B(N531), 
        .Y(N592));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I259_un1_Y_0 (.A(N612), .B(
        N628), .Y(ADD_32x32_fast_I259_un1_Y_0));
    AO1C \state_RNI5VA5I[1]  (.A(un5lt31), .B(next_off_div_2_sqmuxa_11)
        , .C(\state[1]_net_1 ), .Y(un1_state_2_0));
    DFN1E0C0 \off_div[3]  (.D(\next_off_div[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[3]));
    OA1 \off_div_RNI4BJS1[1]  (.A(un5lto4), .B(un5lt4), .C(un5lto7_1), 
        .Y(un5lt9));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I290_Y (.A(sum_2_0), .B(
        off_div[0]), .C(\un1_sum_adj[0] ), .Y(\un1_off_div_1[0] ));
    XNOR2 un13_nsum_adj_I_56 (.A(sum_19), .B(N_6), .Y(I_56_0));
    MX2 \off_div_RNO[7]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[7] ), .S(\state_d_0[2] ), .Y(\next_off_div[7] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I78_Y (.A(N401), .B(N405), .C(
        N404), .Y(N524));
    DFN1E1C0 \sum_adj[21]  (.D(\nsum_adj_11[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[21]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_3 (.A(N610), .B(N625), 
        .C(ADD_32x32_fast_I258_Y_2), .Y(ADD_32x32_fast_I258_Y_3));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I66_Y (.A(N419), .B(N423), .C(
        N422), .Y(N512));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I270_un1_Y (.A(N634), .B(
        N650), .C(N599), .Y(I270_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I8_G0N (.A(\un1_sum_adj[8] )
        , .B(off_div[8]), .Y(N407));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I224_un1_Y (.A(N624), .B(
        N639), .Y(I224_un1_Y));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I299_Y_0 (.A(off_div[9]), .B(
        \un1_sum_adj[9] ), .Y(ADD_32x32_fast_I299_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I1_G0N (.A(\un1_sum_adj[1] )
        , .B(off_div[1]), .Y(N386));
    XA1 \off_div_RNO[4]  (.A(N663), .B(ADD_32x32_fast_I294_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[4] ));
    DFN1E0C0 \off_div[24]  (.D(\next_off_div[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[24]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I64_Y (.A(N422), .B(N426), .C(
        N425), .Y(N510));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I205_Y (.A(N598), .B(
        \un1_sum_adj[0] ), .C(N597), .Y(N663));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I172_Y (.A(N569), .B(N562), 
        .C(N561), .Y(N627));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I3_G0N (.A(sum_2_0), .B(
        \sum_adj[11]_net_1 ), .C(off_div[3]), .Y(N392));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I134_Y (.A(N522), .B(N519), 
        .C(N518), .Y(N583));
    DFN1E1C0 \sum_adj[16]  (.D(\nsum_adj_11[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[16]_net_1 ));
    NOR3A \off_div_RNIMOK71[30]  (.A(un1_off_divlto31_8), .B(
        off_div[23]), .C(off_div[30]), .Y(un1_off_divlto31_15));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I244_Y (.A(N646), .B(N661), 
        .C(N645), .Y(N787));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I238_un1_Y (.A(N653), .B(
        N638), .Y(I238_un1_Y));
    MX2 \sum_adj_RNO[19]  (.A(sum_19), .B(I_56_0), .S(sum_1_0), .Y(
        \nsum_adj_11[19] ));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y_1 (.A(N488), .B(N484), 
        .C(N557), .Y(ADD_32x32_fast_I261_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I126_Y (.A(N514), .B(N511), 
        .C(N510), .Y(N575));
    NOR3 un13_nsum_adj_I_60 (.A(sum_20), .B(sum_19), .C(sum_18), .Y(
        \DWACT_FINC_E[15] ));
    XA1 \off_div_RNO[30]  (.A(N751), .B(ADD_32x32_fast_I320_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[30] ));
    
endmodule


module integral_calc_13s_4_0(
       avg_old,
       avg_new,
       LED_15_0,
       LED_12_0,
       LED_c_2,
       LED_c_0,
       LED_5_0,
       LED_FB_2,
       LED_FB_0,
       choose,
       choose_0_0,
       average,
       LED_33,
       LED_33_i_0,
       calc_avg,
       avg_done,
       choose_n0,
       dec_constd,
       N_45,
       choose_n1,
       inc_constd,
       choose_n2,
       n_rst_c,
       clk_c
    );
input  [11:0] avg_old;
input  [11:0] avg_new;
input  LED_15_0;
input  LED_12_0;
output LED_c_2;
output LED_c_0;
input  LED_5_0;
input  LED_FB_2;
input  LED_FB_0;
input  [2:0] choose;
input  choose_0_0;
output [6:2] average;
output [7:0] LED_33;
output LED_33_i_0;
input  calc_avg;
output avg_done;
output choose_n0;
input  dec_constd;
input  N_45;
output choose_n1;
input  inc_constd;
output choose_n2;
input  n_rst_c;
input  clk_c;

    wire \state_1[0]_net_1 , \state_RNITH201[0]_net_1 , 
        \state_0[0]_net_1 , avg_done_0, \state[1]_net_1 , N649, N529, 
        I192_un1_Y, \un1_integ[8] , N658, ADD_26x26_fast_I238_Y_0, 
        \un1_integ[11] , ADD_26x26_fast_I241_Y_0, N535, I195_un1_Y, 
        \un1_next_int[11] , \state_RNIROBR1[1]_net_1 , 
        ADD_26x26_fast_I253_Y_0, \integ[23]_net_1 , \state[0]_net_1 , 
        ADD_26x26_fast_I254_Y_0, \integ[24]_net_1 , 
        ADD_26x26_fast_I255_Y_0, \integ[25]_net_1 , 
        ADD_26x26_fast_I206_Y_2, N506, N521, ADD_26x26_fast_I206_Y_1, 
        N452, N459, ADD_26x26_fast_I206_Y_0, N402, N398, 
        ADD_26x26_fast_I252_Y_0, \integ[22]_net_1 , 
        ADD_26x26_fast_I205_Y_3, N504, N519, ADD_26x26_fast_I205_Y_2, 
        N450, N457, ADD_26x26_fast_I205_Y_1, ADD_26x26_fast_I205_Y_0, 
        N400, ADD_26x26_fast_I204_Y_3, N502, N517, 
        ADD_26x26_fast_I204_Y_2, N448, N455, ADD_26x26_fast_I204_Y_1, 
        ADD_26x26_fast_I204_Y_0, ADD_26x26_fast_I250_Y_0, 
        \integ[20]_net_1 , ADD_26x26_fast_I251_Y_0, \integ[21]_net_1 , 
        ADD_26x26_fast_I249_Y_0, \integ[19]_net_1 , 
        ADD_26x26_fast_I207_Y_2, N508, N523, ADD_26x26_fast_I207_Y_1, 
        N454, N461, ADD_26x26_fast_I207_Y_0, N404, 
        ADD_26x26_fast_I247_Y_0, \integ[17]_net_1 , 
        ADD_26x26_fast_I246_Y_0, \integ[16]_net_1 , 
        ADD_26x26_fast_I248_Y_0, \integ[18]_net_1 , 
        ADD_26x26_fast_I243_Y_0, ADD_26x26_fast_I209_Y_1, 
        ADD_26x26_fast_I209_un1_Y_0, N543, ADD_26x26_fast_I209_Y_0, 
        N465, N458, ADD_26x26_fast_I208_Y_1, 
        ADD_26x26_fast_I208_un1_Y_0, N541, ADD_26x26_fast_I208_Y_0, 
        N463, N456, ADD_26x26_fast_I239_Y_0, \un18_next_int_m[9] , 
        \inf_abs0_m[9] , ADD_26x26_fast_I210_Y_1, 
        ADD_26x26_fast_I210_un1_Y_0, N491, ADD_26x26_fast_I210_Y_0, 
        N467, N460, ADD_26x26_fast_I205_un1_Y_0, N520, 
        ADD_26x26_fast_I204_un1_Y_0, N518, ADD_26x26_fast_I240_Y_0, 
        \un1_next_int[10] , ADD_26x26_fast_I211_Y_1, 
        ADD_26x26_fast_I211_un1_Y_0, N516, ADD_26x26_fast_I211_Y_0, 
        N469, N462, ADD_26x26_fast_I213_Y_0, 
        ADD_26x26_fast_I213_un1_Y_0, ADD_26x26_fast_I212_Y_0, 
        ADD_26x26_fast_I212_un1_Y_0, ADD_26x26_fast_I234_Y_0, 
        \un1_next_int[4] , ADD_26x26_fast_I235_Y_0, 
        \un18_next_int_m[5] , \inf_abs0_m[5] , N510, N526, N512, N528, 
        N476, N484, N514, N480, N488, N442, N482, N490, 
        \un1_next_int[0] , N478, N486, N493, ADD_26x26_fast_I232_Y_0, 
        \un1_next_int[2] , ADD_26x26_fast_I231_Y_0, \inf_abs0_m[1] , 
        \un18_next_int_m[1] , \integ[1]_net_1 , 
        ADD_26x26_fast_I230_Y_0, \integ[0]_net_1 , 
        ADD_26x26_fast_I77_Y_0, ADD_26x26_fast_I79_Y_0, 
        \un1_integ[15] , \integ[15]_net_1 , N637, \un1_integ[7] , 
        \un1_next_int[7] , N537, I205_un1_Y, N401, I206_un1_Y, N522, 
        \un1_integ[23] , \un1_integ[19] , I180_un1_Y, \un1_integ[24] , 
        \un1_integ[14] , N640, \un1_integ[18] , I182_un1_Y, 
        \un1_integ[21] , I176_un1_Y, \un1_integ[22] , I207_un1_Y, 
        \un1_integ[20] , I178_un1_Y, N524, N539, N399, I204_un1_Y, 
        N533, I194_un1_Y, \un1_integ[3] , \state_RNIHEBR1[1]_net_1 , 
        \un1_integ[25] , \un1_integ[17] , I184_un1_Y, \un1_integ[13] , 
        N525, I190_un1_Y, \un1_integ[4] , \un1_integ[6] , 
        \state_RNINKBR1[0]_net_1 , \un1_integ[2] , \un1_integ[16] , 
        I186_un1_Y, \un1_integ[12] , N646, ADD_26x26_fast_I230_Y, 
        \un1_integ[10] , N531, I193_un1_Y, \un1_integ[9] , 
        \un1_integ[5] , \un1_integ[1] , choose_c1, choose_c0, N_61, 
        N_53, N_69, \inf_abs0_m[8] , \inf_abs0_m[4] , 
        \un18_next_int_m[4] , N_59, N_51, N_35, N_43, N_67, N_98, 
        \inf_abs0_m[6] , \un18_next_int_m[6] , N407, N411, N418, N415, 
        N414, I148_un1_Y, N471, N472, N479, N475, N426, N423, N422, 
        N419, N468, N403, N464, \inf_abs0_m[3] , N474, N489, N481, 
        I163_un1_Y, N527, I108_un1_Y, N430, N427, N342, N339, N431, 
        N333, N473, N420, N347, N351, N350, N421, N425, N470, N417, 
        N429, N466, N440, N437, N436, N441, N318, N321, N433, N432, 
        N428, N332, N483, N434, N348, N329, N477, N424, N485, 
        I121_un1_Y, N345, N344, \inf_abs0_m[2] , \un18_next_int_m[2] , 
        \inf_abs0_m[10] , \un18_next_int_m[10] , I154_un1_Y, N317, 
        N320, N327, N323, N326, N438, N435, N439, N487, N357, N410, 
        N409, \inf_abs0_m[0] , \un18_next_int_m[0] , \inf_abs0_m[11] , 
        N354, N353, N406, I162_un1_Y, I74_un1_Y, N405, N413, N408, 
        \state_RNO_1[1] , N412, N335, N338, \inf_abs0_m[7] , 
        \un18_next_int_m[7] , N341, I152_un1_Y, N416, GND, VCC;
    
    AO1 un1_integ_0_0_ADD_26x26_fast_I56_Y (.A(N341), .B(N345), .C(
        N344), .Y(N424));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I148_un1_Y (.A(N472), .B(N479), 
        .Y(I148_un1_Y));
    DFN1C0 \state[0]  (.D(\state_RNITH201[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state[0]_net_1 ));
    AX1D un1_integ_0_0_choose_n0 (.A(inc_constd), .B(dec_constd), .C(
        choose[0]), .Y(choose_n0));
    DFN1E0C0 \integ[13]  (.D(\un1_integ[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_33[6]));
    DFN1E0C0 \integ[24]  (.D(\un1_integ[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[24]_net_1 ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I61_Y (.A(average[6]), .B(
        \state_RNINKBR1[0]_net_1 ), .C(N339), .Y(N429));
    OR2 un1_integ_0_0_ADD_26x26_fast_I7_P0N (.A(\un1_next_int[7] ), .B(
        LED_33[0]), .Y(N339));
    NOR2A \un1_integ_0_0_LED_5[1]  (.A(LED_33[1]), .B(choose[2]), .Y(
        N_59));
    MX2 \un1_integ_0_0_LED_3[1]  (.A(N_98), .B(N_35), .S(choose[1]), 
        .Y(N_43));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I248_Y_0 (.A(\integ[18]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I248_Y_0));
    MX2 \un1_integ_0_0_LED_6[1]  (.A(N_51), .B(N_59), .S(choose[1]), 
        .Y(N_67));
    AO1B un1_integ_0_0_ADD_26x26_fast_I41_Y (.A(\integ[16]_net_1 ), .B(
        \integ[17]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N409));
    NOR2A \state_RNIOS1U[1]  (.A(\state[1]_net_1 ), .B(avg_old[0]), .Y(
        \un18_next_int_m[0] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I204_un1_Y (.A(N533), .B(
        I194_un1_Y), .C(ADD_26x26_fast_I204_un1_Y_0), .Y(I204_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I86_Y (.A(N408), .B(N404), .Y(
        N457));
    AO1 un1_integ_0_0_ADD_26x26_fast_I98_Y (.A(N420), .B(N417), .C(
        N416), .Y(N469));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I176_un1_Y (.A(N525), .B(N510), 
        .Y(I176_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I205_un1_Y_0 (.A(N504), .B(N520)
        , .Y(ADD_26x26_fast_I205_un1_Y_0));
    OR2 \state_RNIDH661[0]  (.A(\un18_next_int_m[10] ), .B(
        \inf_abs0_m[10] ), .Y(\un1_next_int[10] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I51_Y (.A(N354), .B(N351), .Y(
        N419));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y (.A(
        ADD_26x26_fast_I230_Y_0), .B(\un1_next_int[0] ), .Y(
        ADD_26x26_fast_I230_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I253_Y (.A(I206_un1_Y), .B(
        ADD_26x26_fast_I206_Y_2), .C(ADD_26x26_fast_I253_Y_0), .Y(
        \un1_integ[23] ));
    DFN1E0C0 \integ[21]  (.D(\un1_integ[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[21]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I190_un1_Y (.A(N526), .B(N541), 
        .Y(I190_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I146_Y (.A(N477), .B(N470), .C(
        N469), .Y(N523));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I210_un1_Y_0 (.A(N476), .B(N484)
        , .C(N514), .Y(ADD_26x26_fast_I210_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I142_Y (.A(N473), .B(N466), .C(
        N465), .Y(N519));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I231_Y (.A(
        ADD_26x26_fast_I231_Y_0), .B(N442), .Y(\un1_integ[1] ));
    MX2 \un1_integ_0_0_LED_6[3]  (.A(N_53), .B(N_61), .S(choose[1]), 
        .Y(N_69));
    NOR2A \state_RNI162U[1]  (.A(\state[1]_net_1 ), .B(avg_old[9]), .Y(
        \un18_next_int_m[9] ));
    DFN1E0C0 \integ[15]  (.D(\un1_integ[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[15]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I103_Y (.A(N421), .B(N425), .Y(
        N474));
    NOR2B \state_RNIPH9T[0]  (.A(avg_new[6]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[6] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I125_Y (.A(N448), .B(N456), .Y(
        N502));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_1 (.A(
        ADD_26x26_fast_I209_un1_Y_0), .B(N543), .C(
        ADD_26x26_fast_I209_Y_0), .Y(ADD_26x26_fast_I209_Y_1));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I97_Y (.A(N419), .B(N415), .Y(
        N468));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I77_Y (.A(
        ADD_26x26_fast_I77_Y_0), .B(N399), .Y(N448));
    AO1 un1_integ_0_0_ADD_26x26_fast_I94_Y (.A(N416), .B(N413), .C(
        N412), .Y(N465));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I81_Y (.A(N399), .B(N403), .Y(
        N452));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I151_Y (.A(N482), .B(N474), .Y(
        N528));
    OR2 un1_integ_0_0_ADD_26x26_fast_I74_Y (.A(I74_un1_Y), .B(N317), 
        .Y(N442));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I238_Y (.A(N658), .B(
        ADD_26x26_fast_I238_Y_0), .Y(\un1_integ[8] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I121_Y (.A(I121_un1_Y), .B(N440), 
        .Y(N493));
    AO1A \state_RNIFJ661[1]  (.A(avg_old[11]), .B(\state[1]_net_1 ), 
        .C(\inf_abs0_m[11] ), .Y(\un1_next_int[11] ));
    NOR2B \state_RNI5VEM[0]  (.A(avg_new[11]), .B(\state[0]_net_1 ), 
        .Y(\inf_abs0_m[11] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I154_un1_Y (.A(N485), .B(N478), 
        .Y(I154_un1_Y));
    OR3 un1_integ_0_0_ADD_26x26_fast_I5_P0N (.A(\un18_next_int_m[5] ), 
        .B(\inf_abs0_m[5] ), .C(average[5]), .Y(N333));
    NOR2A \state_RNIV32U[1]  (.A(\state[1]_net_1 ), .B(avg_old[7]), .Y(
        \un18_next_int_m[7] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I246_Y (.A(I186_un1_Y), .B(
        ADD_26x26_fast_I213_Y_0), .C(ADD_26x26_fast_I246_Y_0), .Y(
        \un1_integ[16] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I252_Y_0 (.A(\integ[22]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I252_Y_0));
    DFN1C0 \state_1[0]  (.D(\state_RNITH201[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_1[0]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I39_Y (.A(\integ[17]_net_1 ), .B(
        \integ[18]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N407));
    OA1B un1_integ_0_0_ADD_26x26_fast_I32_Y (.A(\integ[20]_net_1 ), .B(
        \integ[21]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N400));
    NOR2A \state_RNIQU1U[1]  (.A(\state[1]_net_1 ), .B(avg_old[2]), .Y(
        \un18_next_int_m[2] ));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I194_un1_Y (.A(N480), .B(N488), 
        .C(N442), .Y(I194_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I108_un1_Y (.A(N430), .B(N427), 
        .Y(I108_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I100_Y (.A(N419), .B(N422), .C(
        N418), .Y(N471));
    OR2 un1_integ_0_0_ADD_26x26_fast_I12_P0N (.A(LED_33[5]), .B(
        \state[1]_net_1 ), .Y(N354));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I10_G0N (.A(\un1_next_int[10] ), 
        .B(LED_33[3]), .Y(N347));
    DFN1E0C0 \integ[12]  (.D(\un1_integ[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_33[5]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I109_Y (.A(N431), .B(N427), .Y(
        N480));
    MX2 \un1_integ_0_0_LED_1[1]  (.A(LED_12_0), .B(LED_15_0), .S(
        choose_0_0), .Y(N_98));
    OA1B un1_integ_0_0_ADD_26x26_fast_I205_Y_0 (.A(\integ[22]_net_1 ), 
        .B(\integ[23]_net_1 ), .C(\state_0[0]_net_1 ), .Y(
        ADD_26x26_fast_I205_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I115_Y (.A(N437), .B(N433), .Y(
        N486));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I12_G0N (.A(LED_33[5]), .B(
        \state[1]_net_1 ), .Y(N353));
    NOR2A \state_RNIT12U[1]  (.A(\state[1]_net_1 ), .B(avg_old[5]), .Y(
        \un18_next_int_m[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_0 (.A(N463), .B(N456), .C(
        N455), .Y(ADD_26x26_fast_I208_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I111_Y (.A(N433), .B(N429), .Y(
        N482));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I250_Y_0 (.A(\integ[20]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I250_Y_0));
    NOR2B \state_RNIQI9T[0]  (.A(avg_new[7]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[7] ));
    DFN1E0C0 \integ[10]  (.D(\un1_integ[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_33[3]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I180_un1_Y (.A(N514), .B(N529), 
        .Y(I180_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I162_Y (.A(I162_un1_Y), .B(N487), 
        .Y(N541));
    NOR2A \un1_integ_0_0_LED_5[3]  (.A(LED_33[3]), .B(choose[2]), .Y(
        N_61));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I6_G0N (.A(
        \state_RNINKBR1[0]_net_1 ), .B(average[6]), .Y(N335));
    AX1D un1_integ_0_0_ADD_26x26_fast_I249_Y (.A(I180_un1_Y), .B(
        ADD_26x26_fast_I210_Y_1), .C(ADD_26x26_fast_I249_Y_0), .Y(
        \un1_integ[19] ));
    GND GND_i (.Y(GND));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I246_Y_0 (.A(\integ[16]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I246_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I212_un1_Y_0 (.A(N480), .B(N488)
        , .C(N442), .Y(ADD_26x26_fast_I212_un1_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I1_G0N (.A(\inf_abs0_m[1] ), .B(
        \un18_next_int_m[1] ), .C(\integ[1]_net_1 ), .Y(N320));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I107_Y (.A(N425), .B(N429), .Y(
        N478));
    OA1B un1_integ_0_0_ADD_26x26_fast_I38_Y (.A(\integ[17]_net_1 ), .B(
        \integ[18]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N406));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I209_un1_Y_0 (.A(N512), .B(N528)
        , .Y(ADD_26x26_fast_I209_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_3 (.A(N504), .B(N519), .C(
        ADD_26x26_fast_I205_Y_2), .Y(ADD_26x26_fast_I205_Y_3));
    AX1D un1_integ_0_0_ADD_26x26_fast_I255_Y (.A(I204_un1_Y), .B(
        ADD_26x26_fast_I204_Y_3), .C(ADD_26x26_fast_I255_Y_0), .Y(
        \un1_integ[25] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I204_Y_0 (.A(\integ[24]_net_1 ), 
        .B(\integ[23]_net_1 ), .C(\state_1[0]_net_1 ), .Y(
        ADD_26x26_fast_I204_Y_0));
    NOR2B \state_RNIRJ9T[0]  (.A(avg_new[8]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[8] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I243_Y (.A(N525), .B(I190_un1_Y), 
        .C(ADD_26x26_fast_I243_Y_0), .Y(\un1_integ[13] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I231_Y_0 (.A(\inf_abs0_m[1] ), 
        .B(\un18_next_int_m[1] ), .C(\integ[1]_net_1 ), .Y(
        ADD_26x26_fast_I231_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I69_Y (.A(average[2]), .B(
        \un1_next_int[2] ), .C(N327), .Y(N437));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I62_Y (.A(N332), .B(average[6]), 
        .C(\state_RNINKBR1[0]_net_1 ), .Y(N430));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I193_un1_Y (.A(N478), .B(N486), 
        .C(N493), .Y(I193_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I152_un1_Y (.A(N483), .B(N476), 
        .Y(I152_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I7_G0N (.A(\un1_next_int[7] ), 
        .B(LED_33[0]), .Y(N338));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I49_Y (.A(N357), .B(N354), .Y(
        N417));
    OA1B un1_integ_0_0_ADD_26x26_fast_I42_Y (.A(\integ[15]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N410));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I145_Y (.A(N468), .B(N476), .Y(
        N522));
    OR2 un1_integ_0_0_ADD_26x26_fast_I10_P0N (.A(\un1_next_int[10] ), 
        .B(LED_33[3]), .Y(N348));
    OR3 un1_integ_0_0_ADD_26x26_fast_I1_P0N (.A(\inf_abs0_m[1] ), .B(
        \un18_next_int_m[1] ), .C(\integ[1]_net_1 ), .Y(N321));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I184_un1_Y (.A(N533), .B(N518), 
        .Y(I184_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I192_un1_Y (.A(N476), .B(N484), 
        .C(N491), .Y(I192_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I141_Y (.A(N464), .B(N472), .Y(
        N518));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I93_Y (.A(N415), .B(N411), .Y(
        N464));
    AO1B un1_integ_0_0_ADD_26x26_fast_I37_Y (.A(\integ[19]_net_1 ), .B(
        \integ[18]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N405));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I0_G0N (.A(\integ[0]_net_1 ), 
        .B(\state[1]_net_1 ), .Y(N317));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I73_Y (.A(N318), .B(N321), .Y(
        N441));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I59_Y (.A(N342), .B(N339), .Y(
        N427));
    AO1 un1_integ_0_0_ADD_26x26_fast_I52_Y (.A(N347), .B(N351), .C(
        N350), .Y(N420));
    NOR2A \state_RNO[1]  (.A(\state_1[0]_net_1 ), .B(\state[1]_net_1 ), 
        .Y(\state_RNO_1[1] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I34_Y (.A(\integ[19]_net_1 ), .B(
        \integ[20]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N402));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I236_Y (.A(
        \state_RNINKBR1[0]_net_1 ), .B(average[6]), .C(N539), .Y(
        \un1_integ[6] ));
    MX2 \un1_integ_0_0_LED_7[3]  (.A(N_45), .B(N_69), .S(choose[0]), 
        .Y(LED_c_2));
    OR2 un1_integ_0_0_ADD_26x26_fast_I205_Y_1 (.A(
        ADD_26x26_fast_I205_Y_0), .B(N400), .Y(ADD_26x26_fast_I205_Y_1)
        );
    AO1 un1_integ_0_0_ADD_26x26_fast_I150_Y (.A(N481), .B(N474), .C(
        N473), .Y(N527));
    DFN1C0 \integ[0]  (.D(ADD_26x26_fast_I230_Y), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\integ[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I120_Y (.A(N439), .B(N442), .C(
        N438), .Y(N491));
    AO1 un1_integ_0_0_ADD_26x26_fast_I104_Y (.A(N426), .B(N423), .C(
        N422), .Y(N475));
    NOR2B \state_RNILD9T[0]  (.A(avg_new[2]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[2] ));
    VCC VCC_i (.Y(VCC));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I129_Y (.A(N452), .B(N460), .Y(
        N506));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I113_Y (.A(N435), .B(N431), .Y(
        N484));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I241_Y_0 (.A(\un1_next_int[11] ), 
        .B(LED_33[4]), .Y(ADD_26x26_fast_I241_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I89_Y (.A(N407), .B(N411), .Y(
        N460));
    AO1 un1_integ_0_0_ADD_26x26_fast_I68_Y (.A(N323), .B(N327), .C(
        N326), .Y(N436));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_0 (.A(N469), .B(N462), .C(
        N461), .Y(ADD_26x26_fast_I211_Y_0));
    DFN1E0C0 \integ[4]  (.D(\un1_integ[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[4]));
    OR2 un1_integ_0_0_ADD_26x26_fast_I108_Y (.A(I108_un1_Y), .B(N426), 
        .Y(N479));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I3_G0N (.A(
        \state_RNIHEBR1[1]_net_1 ), .B(average[3]), .Y(N326));
    OR2 \state_1_RNIRP8J1[0]  (.A(\un18_next_int_m[0] ), .B(
        \inf_abs0_m[0] ), .Y(\un1_next_int[0] ));
    AO13 un1_integ_0_0_ADD_26x26_fast_I48_Y (.A(LED_33[6]), .B(N353), 
        .C(\state_1[0]_net_1 ), .Y(N416));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I195_un1_Y (.A(N482), .B(N490), 
        .C(\un1_next_int[0] ), .Y(I195_un1_Y));
    DFN1E0C0 \integ[3]  (.D(\un1_integ[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[3]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I252_Y (.A(I207_un1_Y), .B(
        ADD_26x26_fast_I207_Y_2), .C(ADD_26x26_fast_I252_Y_0), .Y(
        \un1_integ[22] ));
    NOR2B \state_RNITH201[0]  (.A(avg_done), .B(calc_avg), .Y(
        \state_RNITH201[0]_net_1 ));
    AO13 un1_integ_0_0_choose_c1 (.A(choose_c0), .B(choose[1]), .C(
        inc_constd), .Y(choose_c1));
    NOR2B \state_1_RNI3T6L[0]  (.A(avg_new[0]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[0] ));
    DFN1E0C0 \integ[6]  (.D(\un1_integ[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[6]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_1 (.A(
        ADD_26x26_fast_I210_un1_Y_0), .B(N491), .C(
        ADD_26x26_fast_I210_Y_0), .Y(ADD_26x26_fast_I210_Y_1));
    AO1A \state_RNIROBR1[1]  (.A(avg_old[8]), .B(\state[1]_net_1 ), .C(
        \inf_abs0_m[8] ), .Y(\state_RNIROBR1[1]_net_1 ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y (.A(N533), .B(I194_un1_Y), 
        .C(ADD_26x26_fast_I239_Y_0), .Y(\un1_integ[9] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I206_Y_0 (.A(N402), .B(N398), .Y(
        ADD_26x26_fast_I206_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I58_Y (.A(N338), .B(N342), .C(
        N341), .Y(N426));
    MX2 \un1_integ_0_0_LED_7[1]  (.A(N_43), .B(N_67), .S(choose[0]), 
        .Y(LED_c_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I67_Y (.A(average[4]), .B(
        \un1_next_int[4] ), .C(N327), .Y(N435));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I253_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I253_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I64_Y (.A(N329), .B(N333), .C(
        N332), .Y(N432));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I204_un1_Y_0 (.A(N502), .B(N518)
        , .Y(ADD_26x26_fast_I204_un1_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I127_Y (.A(N450), .B(N458), .Y(
        N504));
    AO1 un1_integ_0_0_ADD_26x26_fast_I110_Y (.A(N432), .B(N429), .C(
        N428), .Y(N481));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I211_un1_Y_0 (.A(N478), .B(N486)
        , .C(N493), .Y(ADD_26x26_fast_I211_un1_Y_0));
    NOR2A \state_RNI9JNF[1]  (.A(\state[1]_net_1 ), .B(avg_old[10]), 
        .Y(\un18_next_int_m[10] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I90_Y (.A(N412), .B(N408), .Y(
        N461));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I233_Y (.A(
        \state_RNIHEBR1[1]_net_1 ), .B(average[3]), .C(N491), .Y(
        \un1_integ[3] ));
    OA1A un1_integ_0_0_ADD_26x26_fast_I47_Y (.A(\state_1[0]_net_1 ), 
        .B(LED_33[7]), .C(N357), .Y(N415));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I119_Y (.A(N441), .B(N437), .Y(
        N490));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I70_Y (.A(N320), .B(average[2]), 
        .C(\un1_next_int[2] ), .Y(N438));
    DFN1E0C0 \integ[5]  (.D(\un1_integ[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[5]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I182_un1_Y (.A(N516), .B(N531), 
        .Y(I182_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I161_Y (.A(N486), .B(N493), .C(
        N485), .Y(N539));
    OA1B un1_integ_0_0_ADD_26x26_fast_I44_Y (.A(LED_33[7]), .B(
        \integ[15]_net_1 ), .C(\state_1[0]_net_1 ), .Y(N412));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I245_Y (.A(\state_0[0]_net_1 ), 
        .B(\integ[15]_net_1 ), .C(N637), .Y(\un1_integ[15] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I95_Y (.A(N417), .B(N413), .Y(
        N466));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y_0 (.A(
        \un18_next_int_m[9] ), .B(\inf_abs0_m[9] ), .C(LED_33[2]), .Y(
        ADD_26x26_fast_I239_Y_0));
    DFN1E0C0 \integ[2]  (.D(\un1_integ[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[2]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I135_Y (.A(N466), .B(N458), .Y(
        N512));
    OR2 un1_integ_0_0_ADD_26x26_fast_I88_Y (.A(N406), .B(N410), .Y(
        N459));
    AX1D un1_integ_0_0_ADD_26x26_fast_I247_Y (.A(I184_un1_Y), .B(
        ADD_26x26_fast_I212_Y_0), .C(ADD_26x26_fast_I247_Y_0), .Y(
        \un1_integ[17] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I143_Y (.A(N466), .B(N474), .Y(
        N520));
    NOR2B \state_RNIOG9T[0]  (.A(avg_new[5]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[5] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I57_Y (.A(N342), .B(N345), .Y(
        N425));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I186_un1_Y (.A(N535), .B(N520), 
        .Y(I186_un1_Y));
    DFN1E0C0 \integ[23]  (.D(\un1_integ[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[23]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I8_P0N (.A(
        \state_RNIROBR1[1]_net_1 ), .B(LED_33[1]), .Y(N342));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_2 (.A(N506), .B(N521), .C(
        ADD_26x26_fast_I206_Y_1), .Y(ADD_26x26_fast_I206_Y_2));
    AO1 un1_integ_0_0_ADD_26x26_fast_I54_Y (.A(N344), .B(N348), .C(
        N347), .Y(N422));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I131_Y (.A(N454), .B(N462), .Y(
        N508));
    NOR2A \state_RNIS02U[1]  (.A(\state[1]_net_1 ), .B(avg_old[4]), .Y(
        \un18_next_int_m[4] ));
    XNOR3 un1_integ_0_0_choose_n1 (.A(choose[1]), .B(inc_constd), .C(
        choose_c0), .Y(choose_n1));
    AX1D un1_integ_0_0_ADD_26x26_fast_I254_Y (.A(I205_un1_Y), .B(
        ADD_26x26_fast_I205_Y_3), .C(ADD_26x26_fast_I254_Y_0), .Y(
        \un1_integ[24] ));
    DFN1E0C0 \integ[19]  (.D(\un1_integ[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[19]_net_1 ));
    NOR2 \state_0_RNIUQQL[0]  (.A(\state[1]_net_1 ), .B(
        \state_0[0]_net_1 ), .Y(avg_done_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I117_Y (.A(N439), .B(N435), .Y(
        N488));
    DFN1E0C0 \integ[17]  (.D(\un1_integ[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[17]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I33_Y (.A(\integ[21]_net_1 ), .B(
        \integ[20]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N401));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I255_Y_0 (.A(\integ[25]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I255_Y_0));
    DFN1E0C0 \integ[14]  (.D(\un1_integ[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_33[7]));
    NOR2A \un1_integ_0_0_LED_2[1]  (.A(LED_5_0), .B(choose_0_0), .Y(
        N_35));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I87_Y (.A(N405), .B(N409), .Y(
        N458));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y_0 (.A(average[2]), .B(
        \un1_next_int[2] ), .Y(ADD_26x26_fast_I232_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I84_Y (.A(N403), .B(N406), .C(
        N402), .Y(N455));
    OR2 un1_integ_0_0_ADD_26x26_fast_I154_Y (.A(I154_un1_Y), .B(N477), 
        .Y(N531));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I11_G0N (.A(\un1_next_int[11] ), 
        .B(LED_33[4]), .Y(N350));
    AO1 un1_integ_0_0_ADD_26x26_fast_I140_Y (.A(N471), .B(N464), .C(
        N463), .Y(N517));
    NOR2B \state_RNINF9T[0]  (.A(avg_new[4]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[4] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I149_Y (.A(N480), .B(N472), .Y(
        N526));
    AO1 un1_integ_0_0_ADD_26x26_fast_I158_Y (.A(N489), .B(N482), .C(
        N481), .Y(N535));
    NOR2 \state_RNIFC0V[0]  (.A(\state[1]_net_1 ), .B(\state[0]_net_1 )
        , .Y(avg_done));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I249_Y_0 (.A(\integ[19]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I249_Y_0));
    DFN1E0C0 \integ[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[25]_net_1 ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I247_Y_0 (.A(\integ[17]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I247_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y_0 (.A(\integ[0]_net_1 ), 
        .B(\state[1]_net_1 ), .Y(ADD_26x26_fast_I230_Y_0));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I242_Y (.A(\state[1]_net_1 ), .B(
        LED_33[5]), .C(N646), .Y(\un1_integ[12] ));
    DFN1E0C0 \integ[11]  (.D(\un1_integ[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_33[4]));
    DFN1E0C0 \integ[16]  (.D(\un1_integ[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[16]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_1 (.A(
        ADD_26x26_fast_I211_un1_Y_0), .B(N516), .C(
        ADD_26x26_fast_I211_Y_0), .Y(ADD_26x26_fast_I211_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I189_Y (.A(N524), .B(N539), .C(
        N523), .Y(N640));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I254_Y_0 (.A(\integ[24]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I254_Y_0));
    NOR2A \un1_integ_0_0_LED_4[1]  (.A(LED_FB_0), .B(choose[2]), .Y(
        N_51));
    OR2 un1_integ_0_0_ADD_26x26_fast_I163_Y (.A(I163_un1_Y), .B(N489), 
        .Y(N543));
    AO1 un1_integ_0_0_ADD_26x26_fast_I96_Y (.A(N418), .B(N415), .C(
        N414), .Y(N467));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I207_un1_Y (.A(N524), .B(N508), 
        .C(N539), .Y(I207_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I2_G0N (.A(\un1_next_int[2] ), 
        .B(average[2]), .Y(N323));
    AO1 un1_integ_0_0_ADD_26x26_fast_I114_Y (.A(N436), .B(N433), .C(
        N432), .Y(N485));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I147_Y (.A(N470), .B(N478), .Y(
        N524));
    DFN1E0C0 \integ[9]  (.D(\un1_integ[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(LED_33[2]));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I235_Y (.A(
        ADD_26x26_fast_I235_Y_0), .B(N541), .Y(\un1_integ[5] ));
    NOR2B \state_RNIME9T[0]  (.A(avg_new[3]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[3] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I212_Y_0 (.A(
        ADD_26x26_fast_I212_un1_Y_0), .B(N518), .C(N517), .Y(
        ADD_26x26_fast_I212_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I63_Y (.A(average[6]), .B(
        \state_RNINKBR1[0]_net_1 ), .C(N333), .Y(N431));
    AO1 un1_integ_0_0_ADD_26x26_fast_I118_Y (.A(N440), .B(N437), .C(
        N436), .Y(N489));
    NOR2B \state_1_RNI4U6L[0]  (.A(avg_new[1]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[1] ));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I237_Y (.A(\un1_next_int[7] ), 
        .B(LED_33[0]), .C(N537), .Y(\un1_integ[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I133_Y (.A(N456), .B(N464), .Y(
        N510));
    OA1B un1_integ_0_0_ADD_26x26_fast_I30_Y (.A(\integ[22]_net_1 ), .B(
        \integ[21]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N398));
    NOR2B \state_RNI4UEM[0]  (.A(avg_new[10]), .B(\state[0]_net_1 ), 
        .Y(\inf_abs0_m[10] ));
    DFN1E0C0 \integ[22]  (.D(\un1_integ[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[22]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I43_Y (.A(\integ[16]_net_1 ), .B(
        \integ[15]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N411));
    OR2 un1_integ_0_0_ADD_26x26_fast_I192_Y (.A(N529), .B(I192_un1_Y), 
        .Y(N649));
    DFN1E0C0 \integ[1]  (.D(\un1_integ[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(\integ[1]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I35_Y (.A(\integ[20]_net_1 ), .B(
        \integ[19]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N403));
    DFN1C0 \state_0[0]  (.D(\state_RNITH201[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_0[0]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I204_Y_1 (.A(
        ADD_26x26_fast_I204_Y_0), .B(N398), .Y(ADD_26x26_fast_I204_Y_1)
        );
    NOR2B un1_integ_0_0_ADD_26x26_fast_I53_Y (.A(N351), .B(N348), .Y(
        N421));
    AO1 un1_integ_0_0_ADD_26x26_fast_I160_Y (.A(N484), .B(N491), .C(
        N483), .Y(N537));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I91_Y (.A(N413), .B(N409), .Y(
        N462));
    AO1B un1_integ_0_0_ADD_26x26_fast_I79_Y_0 (.A(\integ[22]_net_1 ), 
        .B(\integ[23]_net_1 ), .C(\state_1[0]_net_1 ), .Y(
        ADD_26x26_fast_I79_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I250_Y (.A(I178_un1_Y), .B(
        ADD_26x26_fast_I209_Y_1), .C(ADD_26x26_fast_I250_Y_0), .Y(
        \un1_integ[20] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I240_Y_0 (.A(LED_33[3]), .B(
        \un1_next_int[10] ), .Y(ADD_26x26_fast_I240_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_0 (.A(N467), .B(N460), .C(
        N459), .Y(ADD_26x26_fast_I210_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I71_Y (.A(average[2]), .B(
        \un1_next_int[2] ), .C(N321), .Y(N439));
    DFN1E0C0 \integ[20]  (.D(\un1_integ[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[20]_net_1 ));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I244_Y (.A(\state_0[0]_net_1 ), 
        .B(LED_33[7]), .C(N640), .Y(\un1_integ[14] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_1 (.A(N454), .B(N461), .C(
        ADD_26x26_fast_I207_Y_0), .Y(ADD_26x26_fast_I207_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I106_Y (.A(N428), .B(N425), .C(
        N424), .Y(N477));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_1 (.A(
        ADD_26x26_fast_I208_un1_Y_0), .B(N541), .C(
        ADD_26x26_fast_I208_Y_0), .Y(ADD_26x26_fast_I208_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I102_Y (.A(N424), .B(N421), .C(
        N420), .Y(N473));
    AX1D un1_integ_0_0_ADD_26x26_fast_I251_Y (.A(I176_un1_Y), .B(
        ADD_26x26_fast_I208_Y_1), .C(ADD_26x26_fast_I251_Y_0), .Y(
        \un1_integ[21] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I121_un1_Y (.A(N441), .B(
        \un1_next_int[0] ), .Y(I121_un1_Y));
    OR2 \state_RNIPMBR1[0]  (.A(\un18_next_int_m[7] ), .B(
        \inf_abs0_m[7] ), .Y(\un1_next_int[7] ));
    DFN1E0C0 \integ[18]  (.D(\un1_integ[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[18]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I144_Y (.A(N475), .B(N468), .C(
        N467), .Y(N521));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I139_Y (.A(N462), .B(N470), .Y(
        N516));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I83_Y (.A(N401), .B(N405), .Y(
        N454));
    XNOR3 un1_integ_0_0_choose_n2 (.A(choose_0_0), .B(inc_constd), .C(
        choose_c1), .Y(choose_n2));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_0 (.A(N465), .B(N458), .C(
        N457), .Y(ADD_26x26_fast_I209_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I207_Y_0 (.A(N404), .B(N400), .Y(
        ADD_26x26_fast_I207_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I148_Y (.A(I148_un1_Y), .B(N471), 
        .Y(N525));
    AO1A \state_RNIHEBR1[1]  (.A(avg_old[3]), .B(\state[1]_net_1 ), .C(
        \inf_abs0_m[3] ), .Y(\state_RNIHEBR1[1]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I60_Y (.A(N335), .B(N339), .C(
        N338), .Y(N428));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y (.A(
        ADD_26x26_fast_I232_Y_0), .B(N493), .Y(\un1_integ[2] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I204_Y_2 (.A(N448), .B(N455), .C(
        ADD_26x26_fast_I204_Y_1), .Y(ADD_26x26_fast_I204_Y_2));
    DFN1C0 \state[1]  (.D(\state_RNO_1[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[1]_net_1 ));
    OR2 \state_RNINKBR1[0]  (.A(\un18_next_int_m[6] ), .B(
        \inf_abs0_m[6] ), .Y(\state_RNINKBR1[0]_net_1 ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I9_G0N (.A(\un18_next_int_m[9] ), 
        .B(\inf_abs0_m[9] ), .C(LED_33[2]), .Y(N344));
    OA1B un1_integ_0_0_ADD_26x26_fast_I40_Y (.A(\integ[17]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N408));
    OA1 un1_integ_0_0_ADD_26x26_fast_I65_Y (.A(average[4]), .B(
        \un1_next_int[4] ), .C(N333), .Y(N433));
    AO1 un1_integ_0_0_ADD_26x26_fast_I188_Y (.A(N522), .B(N537), .C(
        N521), .Y(N637));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I178_un1_Y (.A(N512), .B(N527), 
        .Y(I178_un1_Y));
    AO1B un1_integ_0_0_ADD_26x26_fast_I45_Y (.A(\integ[15]_net_1 ), .B(
        LED_33[7]), .C(\state_1[0]_net_1 ), .Y(N413));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I137_Y (.A(N468), .B(N460), .Y(
        N514));
    OR2 un1_integ_0_0_ADD_26x26_fast_I3_P0N (.A(
        \state_RNIHEBR1[1]_net_1 ), .B(average[3]), .Y(N327));
    NOR2A \state_RNIU22U[1]  (.A(\state[1]_net_1 ), .B(avg_old[6]), .Y(
        \un18_next_int_m[6] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I50_Y (.A(N350), .B(N354), .C(
        N353), .Y(N418));
    AO1 un1_integ_0_0_ADD_26x26_fast_I204_Y_3 (.A(N502), .B(N517), .C(
        ADD_26x26_fast_I204_Y_2), .Y(ADD_26x26_fast_I204_Y_3));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I74_un1_Y (.A(N318), .B(
        \un1_next_int[0] ), .Y(I74_un1_Y));
    OA1B un1_integ_0_0_ADD_26x26_fast_I36_Y (.A(\integ[18]_net_1 ), .B(
        \integ[19]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N404));
    OR2 un1_integ_0_0_ADD_26x26_fast_I0_P0N (.A(\integ[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(N318));
    AO1B un1_integ_0_0_ADD_26x26_fast_I77_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\integ[24]_net_1 ), .C(\state_1[0]_net_1 ), .Y(
        ADD_26x26_fast_I77_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I55_Y (.A(N348), .B(N345), .Y(
        N423));
    OA1 un1_integ_0_0_ADD_26x26_fast_I205_un1_Y (.A(N535), .B(
        I195_un1_Y), .C(ADD_26x26_fast_I205_un1_Y_0), .Y(I205_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I163_un1_Y (.A(N490), .B(
        \un1_next_int[0] ), .Y(I163_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_1 (.A(N452), .B(N459), .C(
        ADD_26x26_fast_I206_Y_0), .Y(ADD_26x26_fast_I206_Y_1));
    OA1 un1_integ_0_0_ADD_26x26_fast_I5_G0N (.A(\un18_next_int_m[5] ), 
        .B(\inf_abs0_m[5] ), .C(average[5]), .Y(N332));
    NOR2B \state_RNISK9T[0]  (.A(avg_new[9]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[9] ));
    DFN1E0C0 \integ[7]  (.D(\un1_integ[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(LED_33[0]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_2 (.A(N508), .B(N523), .C(
        ADD_26x26_fast_I207_Y_1), .Y(ADD_26x26_fast_I207_Y_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I4_G0N (.A(\un1_next_int[4] ), 
        .B(average[4]), .Y(N329));
    OR2 un1_integ_0_0_ADD_26x26_fast_I195_Y (.A(N535), .B(I195_un1_Y), 
        .Y(N658));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y (.A(
        ADD_26x26_fast_I234_Y_0), .B(N543), .Y(\un1_integ[4] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_2 (.A(N450), .B(N457), .C(
        ADD_26x26_fast_I205_Y_1), .Y(ADD_26x26_fast_I205_Y_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I162_un1_Y (.A(N488), .B(N442), 
        .Y(I162_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I240_Y (.A(N531), .B(I193_un1_Y), 
        .C(ADD_26x26_fast_I240_Y_0), .Y(\un1_integ[10] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I156_Y (.A(N487), .B(N480), .C(
        N479), .Y(N533));
    DFN1E0C0 \integ[8]  (.D(\un1_integ[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(LED_33[1]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I85_Y (.A(N407), .B(N403), .Y(
        N456));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I251_Y_0 (.A(\integ[21]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I251_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I152_Y (.A(I152_un1_Y), .B(N475), 
        .Y(N529));
    OR3 un1_integ_0_0_ADD_26x26_fast_I9_P0N (.A(\un18_next_int_m[9] ), 
        .B(\inf_abs0_m[9] ), .C(LED_33[2]), .Y(N345));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I208_un1_Y_0 (.A(N510), .B(N526)
        , .Y(ADD_26x26_fast_I208_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I191_Y (.A(N528), .B(N543), .C(
        N527), .Y(N646));
    AO1D un1_integ_0_0_choose_c0 (.A(dec_constd), .B(inc_constd), .C(
        choose[0]), .Y(choose_c0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I31_Y (.A(\integ[22]_net_1 ), .B(
        \integ[21]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N399));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I206_un1_Y (.A(N522), .B(N506), 
        .C(N537), .Y(I206_un1_Y));
    NOR2A \state_RNIPT1U[1]  (.A(\state[1]_net_1 ), .B(avg_old[1]), .Y(
        \un18_next_int_m[1] ));
    OR2 \state_RNIJGBR1[0]  (.A(\un18_next_int_m[4] ), .B(
        \inf_abs0_m[4] ), .Y(\un1_next_int[4] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I235_Y_0 (.A(
        \un18_next_int_m[5] ), .B(\inf_abs0_m[5] ), .C(average[5]), .Y(
        ADD_26x26_fast_I235_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I241_Y (.A(N649), .B(
        ADD_26x26_fast_I241_Y_0), .Y(\un1_integ[11] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I11_P0N (.A(\un1_next_int[11] ), 
        .B(LED_33[4]), .Y(N351));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I243_Y_0 (.A(LED_33[6]), .B(
        \state_1[0]_net_1 ), .Y(ADD_26x26_fast_I243_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I105_Y (.A(N423), .B(N427), .Y(
        N476));
    AO1 un1_integ_0_0_ADD_26x26_fast_I213_Y_0 (.A(
        ADD_26x26_fast_I213_un1_Y_0), .B(N520), .C(N519), .Y(
        ADD_26x26_fast_I213_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I238_Y_0 (.A(
        \state_RNIROBR1[1]_net_1 ), .B(LED_33[1]), .Y(
        ADD_26x26_fast_I238_Y_0));
    INV \integ_RNI0AG3[12]  (.A(LED_33[5]), .Y(LED_33_i_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I101_Y (.A(N419), .B(N423), .Y(
        N472));
    OR2 \state_RNIFCBR1[0]  (.A(\un18_next_int_m[2] ), .B(
        \inf_abs0_m[2] ), .Y(\un1_next_int[2] ));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I66_Y (.A(N326), .B(average[4]), 
        .C(\un1_next_int[4] ), .Y(N434));
    AX1D un1_integ_0_0_ADD_26x26_fast_I248_Y (.A(I182_un1_Y), .B(
        ADD_26x26_fast_I211_Y_1), .C(ADD_26x26_fast_I248_Y_0), .Y(
        \un1_integ[18] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I99_Y (.A(N417), .B(N421), .Y(
        N470));
    AO1 un1_integ_0_0_ADD_26x26_fast_I92_Y (.A(N414), .B(N411), .C(
        N410), .Y(N463));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I79_Y (.A(
        ADD_26x26_fast_I79_Y_0), .B(N401), .Y(N450));
    AO1 un1_integ_0_0_ADD_26x26_fast_I72_Y (.A(N317), .B(N321), .C(
        N320), .Y(N440));
    OR2A un1_integ_0_0_ADD_26x26_fast_I13_P0N (.A(\state[0]_net_1 ), 
        .B(LED_33[6]), .Y(N357));
    OA1B un1_integ_0_0_ADD_26x26_fast_I46_Y (.A(LED_33[6]), .B(
        LED_33[7]), .C(\state_1[0]_net_1 ), .Y(N414));
    AO1 un1_integ_0_0_ADD_26x26_fast_I116_Y (.A(N438), .B(N435), .C(
        N434), .Y(N487));
    NOR2A \un1_integ_0_0_LED_4[3]  (.A(LED_FB_2), .B(choose[2]), .Y(
        N_53));
    AO1 un1_integ_0_0_ADD_26x26_fast_I112_Y (.A(N434), .B(N431), .C(
        N430), .Y(N483));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I8_G0N (.A(
        \state_RNIROBR1[1]_net_1 ), .B(LED_33[1]), .Y(N341));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I213_un1_Y_0 (.A(N482), .B(N490)
        , .C(\un1_next_int[0] ), .Y(ADD_26x26_fast_I213_un1_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y_0 (.A(average[4]), .B(
        \un1_next_int[4] ), .Y(ADD_26x26_fast_I234_Y_0));
    
endmodule


module error_sr_13s_5s_0(
       cur_vd,
       avg_new,
       avg_old,
       avg_enable_1,
       avg_enable_0,
       avg_enable,
       n_rst_c,
       clk_c
    );
input  [11:0] cur_vd;
output [11:0] avg_new;
output [11:0] avg_old;
input  avg_enable_1;
input  avg_enable_0;
input  avg_enable;
input  n_rst_c;
input  clk_c;

    wire \sr_3_[0]_net_1 , \sr_3_[1]_net_1 , \sr_3_[2]_net_1 , 
        \sr_3_[3]_net_1 , \sr_3_[4]_net_1 , \sr_3_[5]_net_1 , 
        \sr_3_[6]_net_1 , \sr_3_[7]_net_1 , \sr_3_[8]_net_1 , 
        \sr_3_[9]_net_1 , \sr_3_[10]_net_1 , \sr_3_[11]_net_1 , 
        \sr_2_[0]_net_1 , \sr_2_[1]_net_1 , \sr_2_[2]_net_1 , 
        \sr_2_[3]_net_1 , \sr_2_[4]_net_1 , \sr_2_[5]_net_1 , 
        \sr_2_[6]_net_1 , \sr_2_[7]_net_1 , \sr_2_[8]_net_1 , 
        \sr_2_[9]_net_1 , \sr_2_[10]_net_1 , \sr_2_[11]_net_1 , 
        \sr_1_[0]_net_1 , \sr_1_[1]_net_1 , \sr_1_[2]_net_1 , 
        \sr_1_[3]_net_1 , \sr_1_[4]_net_1 , \sr_1_[5]_net_1 , 
        \sr_1_[6]_net_1 , \sr_1_[7]_net_1 , \sr_1_[8]_net_1 , 
        \sr_1_[9]_net_1 , \sr_1_[10]_net_1 , \sr_1_[11]_net_1 , GND, 
        VCC;
    
    DFN1E1C0 \sr_1_[11]  (.D(avg_new[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[11]_net_1 ));
    DFN1E1C0 \sr_3_[3]  (.D(\sr_2_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[3]_net_1 ));
    DFN1E1C0 \sr_4_[4]  (.D(\sr_3_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[4]));
    DFN1E1C0 \sr_0_[10]  (.D(cur_vd[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(avg_new[10]));
    DFN1E1C0 \sr_4_[8]  (.D(\sr_3_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[8]));
    DFN1E1C0 \sr_4_[0]  (.D(\sr_3_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[0]));
    DFN1E1C0 \sr_1_[2]  (.D(avg_new[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[2]_net_1 ));
    DFN1E1C0 \sr_0_[2]  (.D(cur_vd[2]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[2]));
    DFN1E1C0 \sr_2_[2]  (.D(\sr_1_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[2]_net_1 ));
    DFN1E1C0 \sr_0_[11]  (.D(cur_vd[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(avg_new[11]));
    DFN1E1C0 \sr_1_[3]  (.D(avg_new[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[3]_net_1 ));
    DFN1E1C0 \sr_0_[3]  (.D(cur_vd[3]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[3]));
    DFN1E1C0 \sr_1_[10]  (.D(avg_new[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[10]_net_1 ));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \sr_4_[10]  (.D(\sr_3_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[10]));
    DFN1E1C0 \sr_3_[11]  (.D(\sr_2_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_3_[11]_net_1 ));
    DFN1E1C0 \sr_2_[3]  (.D(\sr_1_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[3]_net_1 ));
    DFN1E1C0 \sr_3_[6]  (.D(\sr_2_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[6]_net_1 ));
    DFN1E1C0 \sr_3_[1]  (.D(\sr_2_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[1]_net_1 ));
    DFN1E1C0 \sr_4_[2]  (.D(\sr_3_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[2]));
    DFN1E1C0 \sr_1_[6]  (.D(avg_new[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[6]_net_1 ));
    DFN1E1C0 \sr_4_[3]  (.D(\sr_3_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[3]));
    DFN1E1C0 \sr_0_[6]  (.D(cur_vd[6]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[6]));
    DFN1E1C0 \sr_3_[9]  (.D(\sr_2_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[9]_net_1 ));
    DFN1E1C0 \sr_1_[1]  (.D(avg_new[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[1]_net_1 ));
    DFN1E1C0 \sr_0_[1]  (.D(cur_vd[1]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[1]));
    DFN1E1C0 \sr_2_[6]  (.D(\sr_1_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[6]_net_1 ));
    DFN1E1C0 \sr_2_[1]  (.D(\sr_1_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[1]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1C0 \sr_3_[5]  (.D(\sr_2_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[5]_net_1 ));
    DFN1E1C0 \sr_3_[7]  (.D(\sr_2_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[7]_net_1 ));
    DFN1E1C0 \sr_1_[9]  (.D(avg_new[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[9]_net_1 ));
    DFN1E1C0 \sr_0_[9]  (.D(cur_vd[9]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[9]));
    DFN1E1C0 \sr_2_[11]  (.D(\sr_1_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[11]_net_1 ));
    DFN1E1C0 \sr_4_[6]  (.D(\sr_3_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[6]));
    DFN1E1C0 \sr_2_[9]  (.D(\sr_1_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[9]_net_1 ));
    DFN1E1C0 \sr_4_[11]  (.D(\sr_3_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[11]));
    DFN1E1C0 \sr_4_[1]  (.D(\sr_3_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[1]));
    DFN1E1C0 \sr_3_[4]  (.D(\sr_2_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[4]_net_1 ));
    DFN1E1C0 \sr_1_[5]  (.D(avg_new[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[5]_net_1 ));
    DFN1E1C0 \sr_0_[5]  (.D(cur_vd[5]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[5]));
    DFN1E1C0 \sr_1_[7]  (.D(avg_new[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[7]_net_1 ));
    DFN1E1C0 \sr_0_[7]  (.D(cur_vd[7]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[7]));
    DFN1E1C0 \sr_3_[8]  (.D(\sr_2_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[8]_net_1 ));
    DFN1E1C0 \sr_3_[0]  (.D(\sr_2_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[0]_net_1 ));
    DFN1E1C0 \sr_2_[5]  (.D(\sr_1_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[5]_net_1 ));
    DFN1E1C0 \sr_2_[7]  (.D(\sr_1_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[7]_net_1 ));
    DFN1E1C0 \sr_4_[9]  (.D(\sr_3_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[9]));
    DFN1E1C0 \sr_1_[4]  (.D(avg_new[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[4]_net_1 ));
    DFN1E1C0 \sr_0_[4]  (.D(cur_vd[4]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[4]));
    DFN1E1C0 \sr_1_[8]  (.D(avg_new[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[8]_net_1 ));
    DFN1E1C0 \sr_1_[0]  (.D(avg_new[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[0]_net_1 ));
    DFN1E1C0 \sr_2_[4]  (.D(\sr_1_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[4]_net_1 ));
    DFN1E1C0 \sr_0_[8]  (.D(cur_vd[8]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[8]));
    DFN1E1C0 \sr_0_[0]  (.D(cur_vd[0]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[0]));
    DFN1E1C0 \sr_4_[5]  (.D(\sr_3_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[5]));
    DFN1E1C0 \sr_2_[8]  (.D(\sr_1_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[8]_net_1 ));
    DFN1E1C0 \sr_2_[0]  (.D(\sr_1_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[0]_net_1 ));
    DFN1E1C0 \sr_4_[7]  (.D(\sr_3_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[7]));
    DFN1E1C0 \sr_3_[10]  (.D(\sr_2_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_3_[10]_net_1 ));
    DFN1E1C0 \sr_3_[2]  (.D(\sr_2_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[2]_net_1 ));
    DFN1E1C0 \sr_2_[10]  (.D(\sr_1_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[10]_net_1 ));
    
endmodule


module error_sr_13s_64s_0(
       sr_old,
       sr_new,
       cur_error,
       sr_prev,
       sr_new_0_0,
       sr_new_1_0,
       int_enable,
       n_rst_c,
       clk_c
    );
output [12:0] sr_old;
output [12:0] sr_new;
input  [12:0] cur_error;
output [12:0] sr_prev;
output sr_new_0_0;
output sr_new_1_0;
input  int_enable;
input  n_rst_c;
input  clk_c;

    wire \sr_9_[0]_net_1 , \sr_8_[0]_net_1 , \sr_9_[1]_net_1 , 
        \sr_8_[1]_net_1 , \sr_9_[2]_net_1 , \sr_8_[2]_net_1 , 
        \sr_9_[3]_net_1 , \sr_8_[3]_net_1 , \sr_9_[4]_net_1 , 
        \sr_8_[4]_net_1 , \sr_9_[5]_net_1 , \sr_8_[5]_net_1 , 
        \sr_9_[6]_net_1 , \sr_8_[6]_net_1 , \sr_9_[7]_net_1 , 
        \sr_8_[7]_net_1 , \sr_9_[8]_net_1 , \sr_8_[8]_net_1 , 
        \sr_9_[9]_net_1 , \sr_8_[9]_net_1 , \sr_9_[10]_net_1 , 
        \sr_8_[10]_net_1 , \sr_9_[11]_net_1 , \sr_8_[11]_net_1 , 
        \sr_9_[12]_net_1 , \sr_8_[12]_net_1 , \sr_7_[0]_net_1 , 
        \sr_7_[1]_net_1 , \sr_7_[2]_net_1 , \sr_7_[3]_net_1 , 
        \sr_7_[4]_net_1 , \sr_7_[5]_net_1 , \sr_7_[6]_net_1 , 
        \sr_7_[7]_net_1 , \sr_7_[8]_net_1 , \sr_7_[9]_net_1 , 
        \sr_7_[10]_net_1 , \sr_7_[11]_net_1 , \sr_7_[12]_net_1 , 
        \sr_6_[0]_net_1 , \sr_6_[1]_net_1 , \sr_6_[2]_net_1 , 
        \sr_6_[3]_net_1 , \sr_6_[4]_net_1 , \sr_6_[5]_net_1 , 
        \sr_6_[6]_net_1 , \sr_6_[7]_net_1 , \sr_6_[8]_net_1 , 
        \sr_6_[9]_net_1 , \sr_6_[10]_net_1 , \sr_6_[11]_net_1 , 
        \sr_6_[12]_net_1 , \sr_5_[0]_net_1 , \sr_5_[1]_net_1 , 
        \sr_5_[2]_net_1 , \sr_5_[3]_net_1 , \sr_5_[4]_net_1 , 
        \sr_5_[5]_net_1 , \sr_5_[6]_net_1 , \sr_5_[7]_net_1 , 
        \sr_5_[8]_net_1 , \sr_5_[9]_net_1 , \sr_5_[10]_net_1 , 
        \sr_5_[11]_net_1 , \sr_5_[12]_net_1 , \sr_4_[0]_net_1 , 
        \sr_4_[1]_net_1 , \sr_4_[2]_net_1 , \sr_4_[3]_net_1 , 
        \sr_4_[4]_net_1 , \sr_4_[5]_net_1 , \sr_4_[6]_net_1 , 
        \sr_4_[7]_net_1 , \sr_4_[8]_net_1 , \sr_4_[9]_net_1 , 
        \sr_4_[10]_net_1 , \sr_4_[11]_net_1 , \sr_4_[12]_net_1 , 
        \sr_3_[0]_net_1 , \sr_3_[1]_net_1 , \sr_3_[2]_net_1 , 
        \sr_3_[3]_net_1 , \sr_3_[4]_net_1 , \sr_3_[5]_net_1 , 
        \sr_3_[6]_net_1 , \sr_3_[7]_net_1 , \sr_3_[8]_net_1 , 
        \sr_3_[9]_net_1 , \sr_3_[10]_net_1 , \sr_3_[11]_net_1 , 
        \sr_3_[12]_net_1 , \sr_2_[0]_net_1 , \sr_2_[1]_net_1 , 
        \sr_2_[2]_net_1 , \sr_2_[3]_net_1 , \sr_2_[4]_net_1 , 
        \sr_2_[5]_net_1 , \sr_2_[6]_net_1 , \sr_2_[7]_net_1 , 
        \sr_2_[8]_net_1 , \sr_2_[9]_net_1 , \sr_2_[10]_net_1 , 
        \sr_2_[11]_net_1 , \sr_2_[12]_net_1 , \sr_24_[0]_net_1 , 
        \sr_23_[0]_net_1 , \sr_24_[1]_net_1 , \sr_23_[1]_net_1 , 
        \sr_24_[2]_net_1 , \sr_23_[2]_net_1 , \sr_24_[3]_net_1 , 
        \sr_23_[3]_net_1 , \sr_24_[4]_net_1 , \sr_23_[4]_net_1 , 
        \sr_24_[5]_net_1 , \sr_23_[5]_net_1 , \sr_24_[6]_net_1 , 
        \sr_23_[6]_net_1 , \sr_24_[7]_net_1 , \sr_23_[7]_net_1 , 
        \sr_24_[8]_net_1 , \sr_23_[8]_net_1 , \sr_24_[9]_net_1 , 
        \sr_23_[9]_net_1 , \sr_24_[10]_net_1 , \sr_23_[10]_net_1 , 
        \sr_24_[11]_net_1 , \sr_23_[11]_net_1 , \sr_24_[12]_net_1 , 
        \sr_23_[12]_net_1 , \sr_22_[0]_net_1 , \sr_22_[1]_net_1 , 
        \sr_22_[2]_net_1 , \sr_22_[3]_net_1 , \sr_22_[4]_net_1 , 
        \sr_22_[5]_net_1 , \sr_22_[6]_net_1 , \sr_22_[7]_net_1 , 
        \sr_22_[8]_net_1 , \sr_22_[9]_net_1 , \sr_22_[10]_net_1 , 
        \sr_22_[11]_net_1 , \sr_22_[12]_net_1 , \sr_21_[0]_net_1 , 
        \sr_21_[1]_net_1 , \sr_21_[2]_net_1 , \sr_21_[3]_net_1 , 
        \sr_21_[4]_net_1 , \sr_21_[5]_net_1 , \sr_21_[6]_net_1 , 
        \sr_21_[7]_net_1 , \sr_21_[8]_net_1 , \sr_21_[9]_net_1 , 
        \sr_21_[10]_net_1 , \sr_21_[11]_net_1 , \sr_21_[12]_net_1 , 
        \sr_20_[0]_net_1 , \sr_20_[1]_net_1 , \sr_20_[2]_net_1 , 
        \sr_20_[3]_net_1 , \sr_20_[4]_net_1 , \sr_20_[5]_net_1 , 
        \sr_20_[6]_net_1 , \sr_20_[7]_net_1 , \sr_20_[8]_net_1 , 
        \sr_20_[9]_net_1 , \sr_20_[10]_net_1 , \sr_20_[11]_net_1 , 
        \sr_20_[12]_net_1 , \sr_19_[0]_net_1 , \sr_19_[1]_net_1 , 
        \sr_19_[2]_net_1 , \sr_19_[3]_net_1 , \sr_19_[4]_net_1 , 
        \sr_19_[5]_net_1 , \sr_19_[6]_net_1 , \sr_19_[7]_net_1 , 
        \sr_19_[8]_net_1 , \sr_19_[9]_net_1 , \sr_19_[10]_net_1 , 
        \sr_19_[11]_net_1 , \sr_19_[12]_net_1 , \sr_18_[0]_net_1 , 
        \sr_18_[1]_net_1 , \sr_18_[2]_net_1 , \sr_18_[3]_net_1 , 
        \sr_18_[4]_net_1 , \sr_18_[5]_net_1 , \sr_18_[6]_net_1 , 
        \sr_18_[7]_net_1 , \sr_18_[8]_net_1 , \sr_18_[9]_net_1 , 
        \sr_18_[10]_net_1 , \sr_18_[11]_net_1 , \sr_18_[12]_net_1 , 
        \sr_17_[0]_net_1 , \sr_17_[1]_net_1 , \sr_17_[2]_net_1 , 
        \sr_17_[3]_net_1 , \sr_17_[4]_net_1 , \sr_17_[5]_net_1 , 
        \sr_17_[6]_net_1 , \sr_17_[7]_net_1 , \sr_17_[8]_net_1 , 
        \sr_17_[9]_net_1 , \sr_17_[10]_net_1 , \sr_17_[11]_net_1 , 
        \sr_17_[12]_net_1 , \sr_16_[0]_net_1 , \sr_16_[1]_net_1 , 
        \sr_16_[2]_net_1 , \sr_16_[3]_net_1 , \sr_16_[4]_net_1 , 
        \sr_16_[5]_net_1 , \sr_16_[6]_net_1 , \sr_16_[7]_net_1 , 
        \sr_16_[8]_net_1 , \sr_16_[9]_net_1 , \sr_16_[10]_net_1 , 
        \sr_16_[11]_net_1 , \sr_16_[12]_net_1 , \sr_15_[0]_net_1 , 
        \sr_15_[1]_net_1 , \sr_15_[2]_net_1 , \sr_15_[3]_net_1 , 
        \sr_15_[4]_net_1 , \sr_15_[5]_net_1 , \sr_15_[6]_net_1 , 
        \sr_15_[7]_net_1 , \sr_15_[8]_net_1 , \sr_15_[9]_net_1 , 
        \sr_15_[10]_net_1 , \sr_15_[11]_net_1 , \sr_15_[12]_net_1 , 
        \sr_14_[0]_net_1 , \sr_14_[1]_net_1 , \sr_14_[2]_net_1 , 
        \sr_14_[3]_net_1 , \sr_14_[4]_net_1 , \sr_14_[5]_net_1 , 
        \sr_14_[6]_net_1 , \sr_14_[7]_net_1 , \sr_14_[8]_net_1 , 
        \sr_14_[9]_net_1 , \sr_14_[10]_net_1 , \sr_14_[11]_net_1 , 
        \sr_14_[12]_net_1 , \sr_13_[0]_net_1 , \sr_13_[1]_net_1 , 
        \sr_13_[2]_net_1 , \sr_13_[3]_net_1 , \sr_13_[4]_net_1 , 
        \sr_13_[5]_net_1 , \sr_13_[6]_net_1 , \sr_13_[7]_net_1 , 
        \sr_13_[8]_net_1 , \sr_13_[9]_net_1 , \sr_13_[10]_net_1 , 
        \sr_13_[11]_net_1 , \sr_13_[12]_net_1 , \sr_12_[0]_net_1 , 
        \sr_12_[1]_net_1 , \sr_12_[2]_net_1 , \sr_12_[3]_net_1 , 
        \sr_12_[4]_net_1 , \sr_12_[5]_net_1 , \sr_12_[6]_net_1 , 
        \sr_12_[7]_net_1 , \sr_12_[8]_net_1 , \sr_12_[9]_net_1 , 
        \sr_12_[10]_net_1 , \sr_12_[11]_net_1 , \sr_12_[12]_net_1 , 
        \sr_11_[0]_net_1 , \sr_11_[1]_net_1 , \sr_11_[2]_net_1 , 
        \sr_11_[3]_net_1 , \sr_11_[4]_net_1 , \sr_11_[5]_net_1 , 
        \sr_11_[6]_net_1 , \sr_11_[7]_net_1 , \sr_11_[8]_net_1 , 
        \sr_11_[9]_net_1 , \sr_11_[10]_net_1 , \sr_11_[11]_net_1 , 
        \sr_11_[12]_net_1 , \sr_10_[0]_net_1 , \sr_10_[1]_net_1 , 
        \sr_10_[2]_net_1 , \sr_10_[3]_net_1 , \sr_10_[4]_net_1 , 
        \sr_10_[5]_net_1 , \sr_10_[6]_net_1 , \sr_10_[7]_net_1 , 
        \sr_10_[8]_net_1 , \sr_10_[9]_net_1 , \sr_10_[10]_net_1 , 
        \sr_10_[11]_net_1 , \sr_10_[12]_net_1 , \sr_39_[0]_net_1 , 
        \sr_38_[0]_net_1 , \sr_39_[1]_net_1 , \sr_38_[1]_net_1 , 
        \sr_39_[2]_net_1 , \sr_38_[2]_net_1 , \sr_39_[3]_net_1 , 
        \sr_38_[3]_net_1 , \sr_39_[4]_net_1 , \sr_38_[4]_net_1 , 
        \sr_39_[5]_net_1 , \sr_38_[5]_net_1 , \sr_39_[6]_net_1 , 
        \sr_38_[6]_net_1 , \sr_39_[7]_net_1 , \sr_38_[7]_net_1 , 
        \sr_39_[8]_net_1 , \sr_38_[8]_net_1 , \sr_39_[9]_net_1 , 
        \sr_38_[9]_net_1 , \sr_39_[10]_net_1 , \sr_38_[10]_net_1 , 
        \sr_39_[11]_net_1 , \sr_38_[11]_net_1 , \sr_39_[12]_net_1 , 
        \sr_38_[12]_net_1 , \sr_37_[0]_net_1 , \sr_37_[1]_net_1 , 
        \sr_37_[2]_net_1 , \sr_37_[3]_net_1 , \sr_37_[4]_net_1 , 
        \sr_37_[5]_net_1 , \sr_37_[6]_net_1 , \sr_37_[7]_net_1 , 
        \sr_37_[8]_net_1 , \sr_37_[9]_net_1 , \sr_37_[10]_net_1 , 
        \sr_37_[11]_net_1 , \sr_37_[12]_net_1 , \sr_36_[0]_net_1 , 
        \sr_36_[1]_net_1 , \sr_36_[2]_net_1 , \sr_36_[3]_net_1 , 
        \sr_36_[4]_net_1 , \sr_36_[5]_net_1 , \sr_36_[6]_net_1 , 
        \sr_36_[7]_net_1 , \sr_36_[8]_net_1 , \sr_36_[9]_net_1 , 
        \sr_36_[10]_net_1 , \sr_36_[11]_net_1 , \sr_36_[12]_net_1 , 
        \sr_35_[0]_net_1 , \sr_35_[1]_net_1 , \sr_35_[2]_net_1 , 
        \sr_35_[3]_net_1 , \sr_35_[4]_net_1 , \sr_35_[5]_net_1 , 
        \sr_35_[6]_net_1 , \sr_35_[7]_net_1 , \sr_35_[8]_net_1 , 
        \sr_35_[9]_net_1 , \sr_35_[10]_net_1 , \sr_35_[11]_net_1 , 
        \sr_35_[12]_net_1 , \sr_34_[0]_net_1 , \sr_34_[1]_net_1 , 
        \sr_34_[2]_net_1 , \sr_34_[3]_net_1 , \sr_34_[4]_net_1 , 
        \sr_34_[5]_net_1 , \sr_34_[6]_net_1 , \sr_34_[7]_net_1 , 
        \sr_34_[8]_net_1 , \sr_34_[9]_net_1 , \sr_34_[10]_net_1 , 
        \sr_34_[11]_net_1 , \sr_34_[12]_net_1 , \sr_33_[0]_net_1 , 
        \sr_33_[1]_net_1 , \sr_33_[2]_net_1 , \sr_33_[3]_net_1 , 
        \sr_33_[4]_net_1 , \sr_33_[5]_net_1 , \sr_33_[6]_net_1 , 
        \sr_33_[7]_net_1 , \sr_33_[8]_net_1 , \sr_33_[9]_net_1 , 
        \sr_33_[10]_net_1 , \sr_33_[11]_net_1 , \sr_33_[12]_net_1 , 
        \sr_32_[0]_net_1 , \sr_32_[1]_net_1 , \sr_32_[2]_net_1 , 
        \sr_32_[3]_net_1 , \sr_32_[4]_net_1 , \sr_32_[5]_net_1 , 
        \sr_32_[6]_net_1 , \sr_32_[7]_net_1 , \sr_32_[8]_net_1 , 
        \sr_32_[9]_net_1 , \sr_32_[10]_net_1 , \sr_32_[11]_net_1 , 
        \sr_32_[12]_net_1 , \sr_31_[0]_net_1 , \sr_31_[1]_net_1 , 
        \sr_31_[2]_net_1 , \sr_31_[3]_net_1 , \sr_31_[4]_net_1 , 
        \sr_31_[5]_net_1 , \sr_31_[6]_net_1 , \sr_31_[7]_net_1 , 
        \sr_31_[8]_net_1 , \sr_31_[9]_net_1 , \sr_31_[10]_net_1 , 
        \sr_31_[11]_net_1 , \sr_31_[12]_net_1 , \sr_30_[0]_net_1 , 
        \sr_30_[1]_net_1 , \sr_30_[2]_net_1 , \sr_30_[3]_net_1 , 
        \sr_30_[4]_net_1 , \sr_30_[5]_net_1 , \sr_30_[6]_net_1 , 
        \sr_30_[7]_net_1 , \sr_30_[8]_net_1 , \sr_30_[9]_net_1 , 
        \sr_30_[10]_net_1 , \sr_30_[11]_net_1 , \sr_30_[12]_net_1 , 
        \sr_29_[0]_net_1 , \sr_29_[1]_net_1 , \sr_29_[2]_net_1 , 
        \sr_29_[3]_net_1 , \sr_29_[4]_net_1 , \sr_29_[5]_net_1 , 
        \sr_29_[6]_net_1 , \sr_29_[7]_net_1 , \sr_29_[8]_net_1 , 
        \sr_29_[9]_net_1 , \sr_29_[10]_net_1 , \sr_29_[11]_net_1 , 
        \sr_29_[12]_net_1 , \sr_28_[0]_net_1 , \sr_28_[1]_net_1 , 
        \sr_28_[2]_net_1 , \sr_28_[3]_net_1 , \sr_28_[4]_net_1 , 
        \sr_28_[5]_net_1 , \sr_28_[6]_net_1 , \sr_28_[7]_net_1 , 
        \sr_28_[8]_net_1 , \sr_28_[9]_net_1 , \sr_28_[10]_net_1 , 
        \sr_28_[11]_net_1 , \sr_28_[12]_net_1 , \sr_27_[0]_net_1 , 
        \sr_27_[1]_net_1 , \sr_27_[2]_net_1 , \sr_27_[3]_net_1 , 
        \sr_27_[4]_net_1 , \sr_27_[5]_net_1 , \sr_27_[6]_net_1 , 
        \sr_27_[7]_net_1 , \sr_27_[8]_net_1 , \sr_27_[9]_net_1 , 
        \sr_27_[10]_net_1 , \sr_27_[11]_net_1 , \sr_27_[12]_net_1 , 
        \sr_26_[0]_net_1 , \sr_26_[1]_net_1 , \sr_26_[2]_net_1 , 
        \sr_26_[3]_net_1 , \sr_26_[4]_net_1 , \sr_26_[5]_net_1 , 
        \sr_26_[6]_net_1 , \sr_26_[7]_net_1 , \sr_26_[8]_net_1 , 
        \sr_26_[9]_net_1 , \sr_26_[10]_net_1 , \sr_26_[11]_net_1 , 
        \sr_26_[12]_net_1 , \sr_25_[0]_net_1 , \sr_25_[1]_net_1 , 
        \sr_25_[2]_net_1 , \sr_25_[3]_net_1 , \sr_25_[4]_net_1 , 
        \sr_25_[5]_net_1 , \sr_25_[6]_net_1 , \sr_25_[7]_net_1 , 
        \sr_25_[8]_net_1 , \sr_25_[9]_net_1 , \sr_25_[10]_net_1 , 
        \sr_25_[11]_net_1 , \sr_25_[12]_net_1 , \sr_54_[0]_net_1 , 
        \sr_53_[0]_net_1 , \sr_54_[1]_net_1 , \sr_53_[1]_net_1 , 
        \sr_54_[2]_net_1 , \sr_53_[2]_net_1 , \sr_54_[3]_net_1 , 
        \sr_53_[3]_net_1 , \sr_54_[4]_net_1 , \sr_53_[4]_net_1 , 
        \sr_54_[5]_net_1 , \sr_53_[5]_net_1 , \sr_54_[6]_net_1 , 
        \sr_53_[6]_net_1 , \sr_54_[7]_net_1 , \sr_53_[7]_net_1 , 
        \sr_54_[8]_net_1 , \sr_53_[8]_net_1 , \sr_54_[9]_net_1 , 
        \sr_53_[9]_net_1 , \sr_54_[10]_net_1 , \sr_53_[10]_net_1 , 
        \sr_54_[11]_net_1 , \sr_53_[11]_net_1 , \sr_54_[12]_net_1 , 
        \sr_53_[12]_net_1 , \sr_52_[0]_net_1 , \sr_52_[1]_net_1 , 
        \sr_52_[2]_net_1 , \sr_52_[3]_net_1 , \sr_52_[4]_net_1 , 
        \sr_52_[5]_net_1 , \sr_52_[6]_net_1 , \sr_52_[7]_net_1 , 
        \sr_52_[8]_net_1 , \sr_52_[9]_net_1 , \sr_52_[10]_net_1 , 
        \sr_52_[11]_net_1 , \sr_52_[12]_net_1 , \sr_51_[0]_net_1 , 
        \sr_51_[1]_net_1 , \sr_51_[2]_net_1 , \sr_51_[3]_net_1 , 
        \sr_51_[4]_net_1 , \sr_51_[5]_net_1 , \sr_51_[6]_net_1 , 
        \sr_51_[7]_net_1 , \sr_51_[8]_net_1 , \sr_51_[9]_net_1 , 
        \sr_51_[10]_net_1 , \sr_51_[11]_net_1 , \sr_51_[12]_net_1 , 
        \sr_50_[0]_net_1 , \sr_50_[1]_net_1 , \sr_50_[2]_net_1 , 
        \sr_50_[3]_net_1 , \sr_50_[4]_net_1 , \sr_50_[5]_net_1 , 
        \sr_50_[6]_net_1 , \sr_50_[7]_net_1 , \sr_50_[8]_net_1 , 
        \sr_50_[9]_net_1 , \sr_50_[10]_net_1 , \sr_50_[11]_net_1 , 
        \sr_50_[12]_net_1 , \sr_49_[0]_net_1 , \sr_49_[1]_net_1 , 
        \sr_49_[2]_net_1 , \sr_49_[3]_net_1 , \sr_49_[4]_net_1 , 
        \sr_49_[5]_net_1 , \sr_49_[6]_net_1 , \sr_49_[7]_net_1 , 
        \sr_49_[8]_net_1 , \sr_49_[9]_net_1 , \sr_49_[10]_net_1 , 
        \sr_49_[11]_net_1 , \sr_49_[12]_net_1 , \sr_48_[0]_net_1 , 
        \sr_48_[1]_net_1 , \sr_48_[2]_net_1 , \sr_48_[3]_net_1 , 
        \sr_48_[4]_net_1 , \sr_48_[5]_net_1 , \sr_48_[6]_net_1 , 
        \sr_48_[7]_net_1 , \sr_48_[8]_net_1 , \sr_48_[9]_net_1 , 
        \sr_48_[10]_net_1 , \sr_48_[11]_net_1 , \sr_48_[12]_net_1 , 
        \sr_47_[0]_net_1 , \sr_47_[1]_net_1 , \sr_47_[2]_net_1 , 
        \sr_47_[3]_net_1 , \sr_47_[4]_net_1 , \sr_47_[5]_net_1 , 
        \sr_47_[6]_net_1 , \sr_47_[7]_net_1 , \sr_47_[8]_net_1 , 
        \sr_47_[9]_net_1 , \sr_47_[10]_net_1 , \sr_47_[11]_net_1 , 
        \sr_47_[12]_net_1 , \sr_46_[0]_net_1 , \sr_46_[1]_net_1 , 
        \sr_46_[2]_net_1 , \sr_46_[3]_net_1 , \sr_46_[4]_net_1 , 
        \sr_46_[5]_net_1 , \sr_46_[6]_net_1 , \sr_46_[7]_net_1 , 
        \sr_46_[8]_net_1 , \sr_46_[9]_net_1 , \sr_46_[10]_net_1 , 
        \sr_46_[11]_net_1 , \sr_46_[12]_net_1 , \sr_45_[0]_net_1 , 
        \sr_45_[1]_net_1 , \sr_45_[2]_net_1 , \sr_45_[3]_net_1 , 
        \sr_45_[4]_net_1 , \sr_45_[5]_net_1 , \sr_45_[6]_net_1 , 
        \sr_45_[7]_net_1 , \sr_45_[8]_net_1 , \sr_45_[9]_net_1 , 
        \sr_45_[10]_net_1 , \sr_45_[11]_net_1 , \sr_45_[12]_net_1 , 
        \sr_44_[0]_net_1 , \sr_44_[1]_net_1 , \sr_44_[2]_net_1 , 
        \sr_44_[3]_net_1 , \sr_44_[4]_net_1 , \sr_44_[5]_net_1 , 
        \sr_44_[6]_net_1 , \sr_44_[7]_net_1 , \sr_44_[8]_net_1 , 
        \sr_44_[9]_net_1 , \sr_44_[10]_net_1 , \sr_44_[11]_net_1 , 
        \sr_44_[12]_net_1 , \sr_43_[0]_net_1 , \sr_43_[1]_net_1 , 
        \sr_43_[2]_net_1 , \sr_43_[3]_net_1 , \sr_43_[4]_net_1 , 
        \sr_43_[5]_net_1 , \sr_43_[6]_net_1 , \sr_43_[7]_net_1 , 
        \sr_43_[8]_net_1 , \sr_43_[9]_net_1 , \sr_43_[10]_net_1 , 
        \sr_43_[11]_net_1 , \sr_43_[12]_net_1 , \sr_42_[0]_net_1 , 
        \sr_42_[1]_net_1 , \sr_42_[2]_net_1 , \sr_42_[3]_net_1 , 
        \sr_42_[4]_net_1 , \sr_42_[5]_net_1 , \sr_42_[6]_net_1 , 
        \sr_42_[7]_net_1 , \sr_42_[8]_net_1 , \sr_42_[9]_net_1 , 
        \sr_42_[10]_net_1 , \sr_42_[11]_net_1 , \sr_42_[12]_net_1 , 
        \sr_41_[0]_net_1 , \sr_41_[1]_net_1 , \sr_41_[2]_net_1 , 
        \sr_41_[3]_net_1 , \sr_41_[4]_net_1 , \sr_41_[5]_net_1 , 
        \sr_41_[6]_net_1 , \sr_41_[7]_net_1 , \sr_41_[8]_net_1 , 
        \sr_41_[9]_net_1 , \sr_41_[10]_net_1 , \sr_41_[11]_net_1 , 
        \sr_41_[12]_net_1 , \sr_40_[0]_net_1 , \sr_40_[1]_net_1 , 
        \sr_40_[2]_net_1 , \sr_40_[3]_net_1 , \sr_40_[4]_net_1 , 
        \sr_40_[5]_net_1 , \sr_40_[6]_net_1 , \sr_40_[7]_net_1 , 
        \sr_40_[8]_net_1 , \sr_40_[9]_net_1 , \sr_40_[10]_net_1 , 
        \sr_40_[11]_net_1 , \sr_40_[12]_net_1 , \sr_62_[0]_net_1 , 
        \sr_62_[1]_net_1 , \sr_62_[2]_net_1 , \sr_62_[3]_net_1 , 
        \sr_62_[4]_net_1 , \sr_62_[5]_net_1 , \sr_62_[6]_net_1 , 
        \sr_62_[7]_net_1 , \sr_62_[8]_net_1 , \sr_62_[9]_net_1 , 
        \sr_62_[10]_net_1 , \sr_62_[11]_net_1 , \sr_62_[12]_net_1 , 
        \sr_61_[0]_net_1 , \sr_61_[1]_net_1 , \sr_61_[2]_net_1 , 
        \sr_61_[3]_net_1 , \sr_61_[4]_net_1 , \sr_61_[5]_net_1 , 
        \sr_61_[6]_net_1 , \sr_61_[7]_net_1 , \sr_61_[8]_net_1 , 
        \sr_61_[9]_net_1 , \sr_61_[10]_net_1 , \sr_61_[11]_net_1 , 
        \sr_61_[12]_net_1 , \sr_60_[0]_net_1 , \sr_60_[1]_net_1 , 
        \sr_60_[2]_net_1 , \sr_60_[3]_net_1 , \sr_60_[4]_net_1 , 
        \sr_60_[5]_net_1 , \sr_60_[6]_net_1 , \sr_60_[7]_net_1 , 
        \sr_60_[8]_net_1 , \sr_60_[9]_net_1 , \sr_60_[10]_net_1 , 
        \sr_60_[11]_net_1 , \sr_60_[12]_net_1 , \sr_59_[0]_net_1 , 
        \sr_59_[1]_net_1 , \sr_59_[2]_net_1 , \sr_59_[3]_net_1 , 
        \sr_59_[4]_net_1 , \sr_59_[5]_net_1 , \sr_59_[6]_net_1 , 
        \sr_59_[7]_net_1 , \sr_59_[8]_net_1 , \sr_59_[9]_net_1 , 
        \sr_59_[10]_net_1 , \sr_59_[11]_net_1 , \sr_59_[12]_net_1 , 
        \sr_58_[0]_net_1 , \sr_58_[1]_net_1 , \sr_58_[2]_net_1 , 
        \sr_58_[3]_net_1 , \sr_58_[4]_net_1 , \sr_58_[5]_net_1 , 
        \sr_58_[6]_net_1 , \sr_58_[7]_net_1 , \sr_58_[8]_net_1 , 
        \sr_58_[9]_net_1 , \sr_58_[10]_net_1 , \sr_58_[11]_net_1 , 
        \sr_58_[12]_net_1 , \sr_57_[0]_net_1 , \sr_57_[1]_net_1 , 
        \sr_57_[2]_net_1 , \sr_57_[3]_net_1 , \sr_57_[4]_net_1 , 
        \sr_57_[5]_net_1 , \sr_57_[6]_net_1 , \sr_57_[7]_net_1 , 
        \sr_57_[8]_net_1 , \sr_57_[9]_net_1 , \sr_57_[10]_net_1 , 
        \sr_57_[11]_net_1 , \sr_57_[12]_net_1 , \sr_56_[0]_net_1 , 
        \sr_56_[1]_net_1 , \sr_56_[2]_net_1 , \sr_56_[3]_net_1 , 
        \sr_56_[4]_net_1 , \sr_56_[5]_net_1 , \sr_56_[6]_net_1 , 
        \sr_56_[7]_net_1 , \sr_56_[8]_net_1 , \sr_56_[9]_net_1 , 
        \sr_56_[10]_net_1 , \sr_56_[11]_net_1 , \sr_56_[12]_net_1 , 
        \sr_55_[0]_net_1 , \sr_55_[1]_net_1 , \sr_55_[2]_net_1 , 
        \sr_55_[3]_net_1 , \sr_55_[4]_net_1 , \sr_55_[5]_net_1 , 
        \sr_55_[6]_net_1 , \sr_55_[7]_net_1 , \sr_55_[8]_net_1 , 
        \sr_55_[9]_net_1 , \sr_55_[10]_net_1 , \sr_55_[11]_net_1 , 
        \sr_55_[12]_net_1 , GND, VCC;
    
    DFN1E1C0 \sr_41_[5]  (.D(\sr_40_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[5]_net_1 ));
    DFN1E1C0 \sr_15_[3]  (.D(\sr_14_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[3]_net_1 ));
    DFN1E1C0 \sr_36_[5]  (.D(\sr_35_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[5]_net_1 ));
    DFN1E1C0 \sr_57_[5]  (.D(\sr_56_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[5]_net_1 ));
    DFN1E1C0 \sr_45_[11]  (.D(\sr_44_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[11]_net_1 ));
    DFN1E1C0 \sr_39_[6]  (.D(\sr_38_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[6]_net_1 ));
    DFN1E1C0 \sr_36_[4]  (.D(\sr_35_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[4]_net_1 ));
    DFN1E1C0 \sr_42_[4]  (.D(\sr_41_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[4]_net_1 ));
    DFN1E1C0 \sr_9_[3]  (.D(\sr_8_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[3]_net_1 ));
    DFN1E1C0 \sr_6_[4]  (.D(\sr_5_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[4]_net_1 ));
    DFN1E1C0 \sr_32_[3]  (.D(\sr_31_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[3]_net_1 ));
    DFN1E1C0 \sr_52_[6]  (.D(\sr_51_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[6]_net_1 ));
    DFN1E1C0 \sr_21_[9]  (.D(\sr_20_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[9]_net_1 ));
    DFN1E1C0 \sr_47_[12]  (.D(\sr_46_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[12]_net_1 ));
    DFN1E1C0 \sr_22_[4]  (.D(\sr_21_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[4]_net_1 ));
    DFN1E1C0 \sr_10_[1]  (.D(\sr_9_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[1]_net_1 ));
    DFN1E1C0 \sr_5_[4]  (.D(\sr_4_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[4]_net_1 ));
    DFN1E1C0 \sr_62_[6]  (.D(\sr_61_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[6]_net_1 ));
    DFN1E1C0 \sr_58_[2]  (.D(\sr_57_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[2]_net_1 ));
    DFN1E1C0 \sr_55_[0]  (.D(\sr_54_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[0]_net_1 ));
    DFN1E1C0 \sr_27_[3]  (.D(\sr_26_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[3]_net_1 ));
    DFN1E1C0 \sr_21_[1]  (.D(\sr_20_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[1]_net_1 ));
    DFN1E1C0 \sr_37_[9]  (.D(\sr_36_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[9]_net_1 ));
    DFN1E1C0 \sr_48_[10]  (.D(\sr_47_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[10]_net_1 ));
    DFN1E1C0 \sr_60_[5]  (.D(\sr_59_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[5]_net_1 ));
    DFN1E1C0 \sr_30_[5]  (.D(\sr_29_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[5]_net_1 ));
    DFN1E1C0 \sr_14_[4]  (.D(\sr_13_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[4]_net_1 ));
    DFN1E1C0 \sr_24_[8]  (.D(\sr_23_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[8]_net_1 ));
    DFN1E1C0 \sr_30_[4]  (.D(\sr_29_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[4]_net_1 ));
    DFN1E1C0 \sr_37_[6]  (.D(\sr_36_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[6]_net_1 ));
    DFN1E1C0 \sr_42_[6]  (.D(\sr_41_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[6]_net_1 ));
    DFN1E1C0 \sr_58_[4]  (.D(\sr_57_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[4]_net_1 ));
    DFN1E1C0 \sr_57_[10]  (.D(\sr_56_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[10]_net_1 ));
    DFN1E1C0 \sr_43_[7]  (.D(\sr_42_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[7]_net_1 ));
    DFN1E1C0 \sr_44_[2]  (.D(\sr_43_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[2]_net_1 ));
    DFN1E1C0 \sr_53_[7]  (.D(\sr_52_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[7]_net_1 ));
    DFN1E1C0 \sr_59_[1]  (.D(\sr_58_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[1]_net_1 ));
    DFN1E1C0 \sr_27_[10]  (.D(\sr_26_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[10]_net_1 ));
    DFN1E1C0 \sr_53_[8]  (.D(\sr_52_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[8]_net_1 ));
    DFN1E1C0 \sr_16_[4]  (.D(\sr_15_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[4]_net_1 ));
    DFN1E1C0 \sr_10_[11]  (.D(\sr_9_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[11]_net_1 ));
    DFN1E1C0 \sr_26_[8]  (.D(\sr_25_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[8]_net_1 ));
    DFN1E1C0 \sr_63_[7]  (.D(\sr_62_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[7]));
    DFN1E1C0 \sr_28_[7]  (.D(\sr_27_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[7]_net_1 ));
    DFN1E1C0 \sr_63_[8]  (.D(\sr_62_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[8]));
    DFN1E1C0 \sr_24_[0]  (.D(\sr_23_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[0]_net_1 ));
    DFN1E1C0 \sr_46_[2]  (.D(\sr_45_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[2]_net_1 ));
    DFN1E1C0 \sr_13_[5]  (.D(\sr_12_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[5]_net_1 ));
    DFN1E1C0 \sr_0_[2]  (.D(cur_error[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[2]));
    DFN1E1C0 \sr_0_[8]  (.D(cur_error[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[8]));
    DFN1E1C0 \sr_8_[3]  (.D(\sr_7_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[3]_net_1 ));
    DFN1E1C0 \sr_42_[11]  (.D(\sr_41_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[11]_net_1 ));
    DFN1E1C0 \sr_13_[3]  (.D(\sr_12_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[3]_net_1 ));
    DFN1E1C0 \sr_54_[10]  (.D(\sr_53_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[10]_net_1 ));
    DFN1E1C0 \sr_37_[11]  (.D(\sr_36_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[11]_net_1 ));
    DFN1E1C0 \sr_19_[7]  (.D(\sr_18_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[7]_net_1 ));
    DFN1E1C0 \sr_57_[1]  (.D(\sr_56_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[1]_net_1 ));
    DFN1E1C0 \sr_44_[11]  (.D(\sr_43_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[11]_net_1 ));
    DFN1E1C0 \sr_32_[10]  (.D(\sr_31_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[10]_net_1 ));
    DFN1E1C0 \sr_26_[0]  (.D(\sr_25_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[0]_net_1 ));
    DFN1E1C0 \sr_24_[10]  (.D(\sr_23_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[10]_net_1 ));
    DFN1E1C0 \sr_12_[1]  (.D(\sr_11_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[1]_net_1 ));
    DFN1E1C0 \sr_10_[4]  (.D(\sr_9_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[4]_net_1 ));
    DFN1E1C0 \sr_63_[0]  (.D(\sr_62_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[0]));
    DFN1E1C0 \sr_20_[8]  (.D(\sr_19_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[8]_net_1 ));
    DFN1E1C0 \sr_60_[12]  (.D(\sr_59_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[12]_net_1 ));
    DFN1E1C0 \sr_6_[10]  (.D(\sr_5_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[10]_net_1 ));
    DFN1E1C0 \sr_19_[6]  (.D(\sr_18_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[6]_net_1 ));
    DFN1E1C0 \sr_62_[5]  (.D(\sr_61_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[5]_net_1 ));
    DFN1E1C0 \sr_44_[8]  (.D(\sr_43_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[8]_net_1 ));
    DFN1E1C0 \sr_49_[5]  (.D(\sr_48_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[5]_net_1 ));
    DFN1E1C0 \sr_53_[0]  (.D(\sr_52_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[0]_net_1 ));
    DFN1E1C0 \sr_1_[2]  (.D(sr_new[2]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[2]));
    DFN1E1C0 \sr_40_[2]  (.D(\sr_39_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[2]_net_1 ));
    DFN1E1C0 \sr_32_[5]  (.D(\sr_31_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[5]_net_1 ));
    DFN1E1C0 \sr_1_[8]  (.D(sr_new[8]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[8]));
    DFN1E1C0 \sr_18_[12]  (.D(\sr_17_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[12]_net_1 ));
    DFN1E1C0 \sr_60_[10]  (.D(\sr_59_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[10]_net_1 ));
    DFN1E1C0 \sr_32_[4]  (.D(\sr_31_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[4]_net_1 ));
    DFN1E1C0 \sr_54_[3]  (.D(\sr_53_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[3]_net_1 ));
    DFN1E1C0 \sr_29_[9]  (.D(\sr_28_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[9]_net_1 ));
    DFN1E1C0 \sr_24_[2]  (.D(\sr_23_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[2]_net_1 ));
    DFN1E1C0 \sr_18_[9]  (.D(\sr_17_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[9]_net_1 ));
    DFN1E1C0 \sr_7_[9]  (.D(\sr_6_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[9]_net_1 ));
    DFN1E1C0 \sr_63_[10]  (.D(\sr_62_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[10]));
    DFN1E1C0 \sr_24_[5]  (.D(\sr_23_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[5]_net_1 ));
    DFN1E1C0 \sr_46_[8]  (.D(\sr_45_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[8]_net_1 ));
    DFN1E1C0 \sr_59_[11]  (.D(\sr_58_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[11]_net_1 ));
    DFN1E1C0 \sr_17_[7]  (.D(\sr_16_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[7]_net_1 ));
    DFN1E1C0 \sr_14_[8]  (.D(\sr_13_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[8]_net_1 ));
    DFN1E1C0 \sr_41_[3]  (.D(\sr_40_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[3]_net_1 ));
    DFN1E1C0 \sr_20_[0]  (.D(\sr_19_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[0]_net_1 ));
    DFN1E1C0 \sr_48_[0]  (.D(\sr_47_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[0]_net_1 ));
    DFN1E1C0 \sr_29_[1]  (.D(\sr_28_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[1]_net_1 ));
    DFN1E1C0 \sr_3_[10]  (.D(\sr_2_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[10]_net_1 ));
    DFN1E1C0 \sr_29_[11]  (.D(\sr_28_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[11]_net_1 ));
    DFN1E1C0 \sr_35_[1]  (.D(\sr_34_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[1]_net_1 ));
    DFN1E1C0 \sr_17_[6]  (.D(\sr_16_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[6]_net_1 ));
    DFN1E1C0 \sr_2_[3]  (.D(sr_prev[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[3]_net_1 ));
    DFN1E1C0 \sr_56_[3]  (.D(\sr_55_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[3]_net_1 ));
    DFN1E1C0 \sr_47_[5]  (.D(\sr_46_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[5]_net_1 ));
    DFN1E1C0 \sr_35_[2]  (.D(\sr_34_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[2]_net_1 ));
    DFN1E1C0 \sr_35_[12]  (.D(\sr_34_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[12]_net_1 ));
    DFN1E1C0 \sr_26_[2]  (.D(\sr_25_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[2]_net_1 ));
    DFN1E1C0 \sr_6_[2]  (.D(\sr_5_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[2]_net_1 ));
    DFN1E1C0 \sr_6_[8]  (.D(\sr_5_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[8]_net_1 ));
    DFN1E1C0 \sr_35_[7]  (.D(\sr_34_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[7]_net_1 ));
    DFN1E1C0 \sr_26_[5]  (.D(\sr_25_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[5]_net_1 ));
    DFN1E1C0 \sr_16_[8]  (.D(\sr_15_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[8]_net_1 ));
    DFN1E1C0 \sr_52_[12]  (.D(\sr_51_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[12]_net_1 ));
    DFN1E1C0 \sr_5_[2]  (.D(\sr_4_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[2]_net_1 ));
    DFN1E1C0 \sr_5_[8]  (.D(\sr_4_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[8]_net_1 ));
    DFN1E1C0 \sr_27_[9]  (.D(\sr_26_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[9]_net_1 ));
    DFN1E1C0 \sr_18_[11]  (.D(\sr_17_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[11]_net_1 ));
    DFN1E1C0 \sr_3_[9]  (.D(\sr_2_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[9]_net_1 ));
    DFN1E1C0 \sr_2_[11]  (.D(sr_prev[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[11]_net_1 ));
    DFN1E1C0 \sr_40_[8]  (.D(\sr_39_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[8]_net_1 ));
    DFN1E1C0 \sr_22_[12]  (.D(\sr_21_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[12]_net_1 ));
    DFN1E1C0 \sr_45_[9]  (.D(\sr_44_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[9]_net_1 ));
    DFN1E1C0 \sr_2_[12]  (.D(sr_prev[12]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[12]_net_1 ));
    DFN1E1C0 \sr_27_[1]  (.D(\sr_26_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[1]_net_1 ));
    DFN1E1C0 \sr_0__1[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_new_1_0));
    DFN1E1C0 \sr_9_[4]  (.D(\sr_8_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[4]_net_1 ));
    DFN1E1C0 \sr_12_[4]  (.D(\sr_11_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[4]_net_1 ));
    DFN1E1C0 \sr_56_[11]  (.D(\sr_55_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[11]_net_1 ));
    DFN1E1C0 \sr_22_[8]  (.D(\sr_21_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[8]_net_1 ));
    DFN1E1C0 \sr_14_[2]  (.D(\sr_13_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[2]_net_1 ));
    DFN1E1C0 \sr_46_[12]  (.D(\sr_45_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[12]_net_1 ));
    DFN1E1C0 \sr_50_[3]  (.D(\sr_49_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[3]_net_1 ));
    DFN1E1C0 \sr_20_[2]  (.D(\sr_19_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[2]_net_1 ));
    DFN1E1C0 \sr_44_[12]  (.D(\sr_43_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[12]_net_1 ));
    DFN1E1C0 \sr_26_[11]  (.D(\sr_25_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[11]_net_1 ));
    DFN1E1C0 \sr_14_[0]  (.D(\sr_13_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[0]_net_1 ));
    DFN1E1C0 \sr_34_[8]  (.D(\sr_33_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[8]_net_1 ));
    DFN1E1C0 \sr_20_[5]  (.D(\sr_19_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[5]_net_1 ));
    DFN1E1C0 \sr_10_[8]  (.D(\sr_9_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[8]_net_1 ));
    DFN1E1C0 \sr_42_[2]  (.D(\sr_41_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[2]_net_1 ));
    DFN1E1C0 \sr_55_[11]  (.D(\sr_54_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[11]_net_1 ));
    DFN1E1C0 \sr_51_[9]  (.D(\sr_50_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[9]_net_1 ));
    DFN1E1C0 \sr_54_[5]  (.D(\sr_53_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[5]_net_1 ));
    DFN1E1C0 \sr_25_[11]  (.D(\sr_24_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[11]_net_1 ));
    DFN1E1C0 \sr_21_[6]  (.D(\sr_20_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[6]_net_1 ));
    DFN1E1C0 \sr_57_[12]  (.D(\sr_56_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[12]_net_1 ));
    DFN1E1C0 \sr_16_[2]  (.D(\sr_15_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[2]_net_1 ));
    DFN1E1C0 \sr_35_[0]  (.D(\sr_34_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[0]_net_1 ));
    DFN1E1C0 \sr_16_[0]  (.D(\sr_15_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[0]_net_1 ));
    DFN1E1C0 \sr_36_[8]  (.D(\sr_35_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[8]_net_1 ));
    DFN1E1C0 \sr_27_[12]  (.D(\sr_26_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[12]_net_1 ));
    DFN1E1C0 \sr_22_[0]  (.D(\sr_21_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[0]_net_1 ));
    DFN1E1C0 \sr_0__0[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_new_0_0));
    DFN1E1C0 \sr_13_[11]  (.D(\sr_12_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[11]_net_1 ));
    DFN1E1C0 \sr_58_[10]  (.D(\sr_57_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[10]_net_1 ));
    DFN1E1C0 \sr_7_[12]  (.D(\sr_6_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[12]_net_1 ));
    DFN1E1C0 \sr_24_[3]  (.D(\sr_23_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[3]_net_1 ));
    DFN1E1C0 \sr_34_[9]  (.D(\sr_33_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[9]_net_1 ));
    DFN1E1C0 \sr_28_[10]  (.D(\sr_27_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[10]_net_1 ));
    DFN1E1C0 \sr_56_[5]  (.D(\sr_55_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[5]_net_1 ));
    DFN1E1C0 \sr_7_[10]  (.D(\sr_6_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[10]_net_1 ));
    DFN1E1C0 \sr_33_[1]  (.D(\sr_32_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[1]_net_1 ));
    DFN1E1C0 \sr_33_[2]  (.D(\sr_32_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[2]_net_1 ));
    DFN1E1C0 \sr_48_[7]  (.D(\sr_47_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[7]_net_1 ));
    DFN1E1C0 \sr_58_[7]  (.D(\sr_57_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[7]_net_1 ));
    DFN1E1C0 \sr_34_[6]  (.D(\sr_33_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[6]_net_1 ));
    DFN1E1C0 \sr_33_[7]  (.D(\sr_32_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[7]_net_1 ));
    DFN1E1C0 \sr_10_[2]  (.D(\sr_9_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[2]_net_1 ));
    DFN1E1C0 \sr_26_[3]  (.D(\sr_25_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[3]_net_1 ));
    DFN1E1C0 \sr_36_[9]  (.D(\sr_35_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[9]_net_1 ));
    DFN1E1C0 \sr_58_[8]  (.D(\sr_57_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[8]_net_1 ));
    DFN1E1C0 \sr_42_[8]  (.D(\sr_41_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[8]_net_1 ));
    DFN1E1C0 \sr_49_[3]  (.D(\sr_48_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[3]_net_1 ));
    DFN1E1C0 \sr_10_[0]  (.D(\sr_9_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[0]_net_1 ));
    DFN1E1C0 \sr_30_[8]  (.D(\sr_29_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[8]_net_1 ));
    DFN1E1C0 \sr_35_[10]  (.D(\sr_34_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[10]_net_1 ));
    DFN1E1C0 \sr_8_[4]  (.D(\sr_7_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[4]_net_1 ));
    DFN1E1C0 \sr_43_[12]  (.D(\sr_42_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[12]_net_1 ));
    DFN1E1C0 \sr_0_[9]  (.D(cur_error[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[9]));
    DFN1E1C0 \sr_43_[9]  (.D(\sr_42_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[9]_net_1 ));
    DFN1E1C0 \sr_50_[5]  (.D(\sr_49_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[5]_net_1 ));
    DFN1E1C0 \sr_52_[3]  (.D(\sr_51_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[3]_net_1 ));
    DFN1E1C0 \sr_22_[2]  (.D(\sr_21_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[2]_net_1 ));
    DFN1E1C0 \sr_18_[5]  (.D(\sr_17_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[5]_net_1 ));
    DFN1E1C0 \sr_7_[0]  (.D(\sr_6_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[0]_net_1 ));
    DFN1E1C0 \sr_36_[6]  (.D(\sr_35_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[6]_net_1 ));
    DFN1E1C0 \sr_60_[11]  (.D(\sr_59_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[11]_net_1 ));
    DFN1E1C0 \sr_45_[4]  (.D(\sr_44_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[4]_net_1 ));
    DFN1E1C0 \sr_22_[5]  (.D(\sr_21_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[5]_net_1 ));
    DFN1E1C0 \sr_35_[3]  (.D(\sr_34_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[3]_net_1 ));
    DFN1E1C0 \sr_7_[6]  (.D(\sr_6_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[6]_net_1 ));
    DFN1E1C0 \sr_12_[8]  (.D(\sr_11_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[8]_net_1 ));
    DFN1E1C0 \sr_55_[6]  (.D(\sr_54_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[6]_net_1 ));
    DFN1E1C0 \sr_52_[11]  (.D(\sr_51_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[11]_net_1 ));
    DFN1E1C0 \sr_18_[3]  (.D(\sr_17_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[3]_net_1 ));
    DFN1E1C0 \sr_36_[10]  (.D(\sr_35_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[10]_net_1 ));
    DFN1E1C0 \sr_25_[4]  (.D(\sr_24_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[4]_net_1 ));
    DFN1E1C0 \sr_22_[11]  (.D(\sr_21_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[11]_net_1 ));
    DFN1E1C0 \sr_20_[3]  (.D(\sr_19_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[3]_net_1 ));
    DFN1E1C0 \sr_30_[9]  (.D(\sr_29_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[9]_net_1 ));
    DFN1E1C0 \sr_47_[3]  (.D(\sr_46_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[3]_net_1 ));
    DFN1E1C0 \sr_54_[11]  (.D(\sr_53_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[11]_net_1 ));
    DFN1E1C0 \sr_4_[7]  (.D(\sr_3_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[7]_net_1 ));
    DFN1E1C0 \sr_31_[12]  (.D(\sr_30_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[12]_net_1 ));
    DFN1E1C0 \sr_54_[1]  (.D(\sr_53_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[1]_net_1 ));
    DFN1E1C0 \sr_24_[11]  (.D(\sr_23_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[11]_net_1 ));
    DFN1E1C0 \sr_1_[9]  (.D(sr_new[9]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[9]));
    DFN1E1C0 \sr_58_[0]  (.D(\sr_57_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[0]_net_1 ));
    DFN1E1C0 \sr_33_[0]  (.D(\sr_32_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[0]_net_1 ));
    DFN1E1C0 \sr_41_[1]  (.D(\sr_40_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[1]_net_1 ));
    DFN1E1C0 \sr_30_[6]  (.D(\sr_29_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[6]_net_1 ));
    DFN1E1C0 \sr_7_[1]  (.D(\sr_6_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[1]_net_1 ));
    DFN1E1C0 \sr_3_[0]  (.D(\sr_2_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[0]_net_1 ));
    DFN1E1C0 \sr_45_[6]  (.D(\sr_44_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[6]_net_1 ));
    DFN1E1C0 \sr_3_[6]  (.D(\sr_2_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[6]_net_1 ));
    DFN1E1C0 \sr_59_[9]  (.D(\sr_58_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[9]_net_1 ));
    DFN1E1C0 \sr_2_[4]  (.D(sr_prev[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[4]_net_1 ));
    DFN1E1C0 \sr_56_[1]  (.D(\sr_55_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[1]_net_1 ));
    DFN1E1C0 \sr_29_[6]  (.D(\sr_28_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[6]_net_1 ));
    DFN1E1C0 \sr_9_[2]  (.D(\sr_8_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[2]_net_1 ));
    DFN1E1C0 \sr_9_[8]  (.D(\sr_8_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[8]_net_1 ));
    DFN1E1C0 \sr_17_[11]  (.D(\sr_16_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[11]_net_1 ));
    DFN1E1C0 \sr_12_[2]  (.D(\sr_11_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[2]_net_1 ));
    DFN1E1C0 \sr_12_[10]  (.D(\sr_11_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[10]_net_1 ));
    DFN1E1C0 \sr_12_[0]  (.D(\sr_11_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[0]_net_1 ));
    DFN1E1C0 \sr_32_[8]  (.D(\sr_31_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[8]_net_1 ));
    DFN1E1C0 \sr_14_[7]  (.D(\sr_13_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[7]_net_1 ));
    DFN1E1C0 \sr_6_[9]  (.D(\sr_5_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[9]_net_1 ));
    DFN1E1C0 \sr_31_[10]  (.D(\sr_30_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[10]_net_1 ));
    DFN1E1C0 \sr_31_[11]  (.D(\sr_30_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[11]_net_1 ));
    DFN1E1C0 \sr_14_[6]  (.D(\sr_13_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[6]_net_1 ));
    DFN1E1C0 \sr_5_[10]  (.D(\sr_4_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[10]_net_1 ));
    DFN1E1C0 \sr_5_[9]  (.D(\sr_4_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[9]_net_1 ));
    DFN1E1C0 \sr_52_[5]  (.D(\sr_51_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[5]_net_1 ));
    DFN1E1C0 \sr_3_[1]  (.D(\sr_2_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[1]_net_1 ));
    DFN1E1C0 \sr_44_[5]  (.D(\sr_43_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[5]_net_1 ));
    DFN1E1C0 \sr_57_[9]  (.D(\sr_56_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[9]_net_1 ));
    DFN1E1C0 \sr_50_[1]  (.D(\sr_49_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[1]_net_1 ));
    DFN1E1C0 \sr_16_[7]  (.D(\sr_15_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[7]_net_1 ));
    DFN1E1C0 \sr_51_[2]  (.D(\sr_50_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[2]_net_1 ));
    DFN1E1C0 \sr_27_[6]  (.D(\sr_26_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[6]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1C0 \sr_43_[4]  (.D(\sr_42_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[4]_net_1 ));
    DFN1E1C0 \sr_24_[9]  (.D(\sr_23_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[9]_net_1 ));
    DFN1E1C0 \sr_22_[3]  (.D(\sr_21_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[3]_net_1 ));
    DFN1E1C0 \sr_33_[3]  (.D(\sr_32_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[3]_net_1 ));
    DFN1E1C0 \sr_32_[9]  (.D(\sr_31_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[9]_net_1 ));
    DFN1E1C0 \sr_15_[1]  (.D(\sr_14_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[1]_net_1 ));
    DFN1E1C0 \sr_53_[6]  (.D(\sr_52_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[6]_net_1 ));
    DFN1E1C0 \sr_60_[1]  (.D(\sr_59_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[1]_net_1 ));
    DFN1E1C0 \sr_16_[6]  (.D(\sr_15_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[6]_net_1 ));
    DFN1E1C0 \sr_61_[2]  (.D(\sr_60_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[2]_net_1 ));
    DFN1E1C0 \sr_23_[4]  (.D(\sr_22_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[4]_net_1 ));
    DFN1E1C0 \sr_46_[5]  (.D(\sr_45_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[5]_net_1 ));
    DFN1E1C0 \sr_24_[1]  (.D(\sr_23_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[1]_net_1 ));
    DFN1E1C0 \sr_63_[6]  (.D(\sr_62_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[6]));
    DFN1E1C0 \sr_49_[12]  (.D(\sr_48_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[12]_net_1 ));
    DFN1E1C0 \sr_56_[12]  (.D(\sr_55_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[12]_net_1 ));
    DFN1E1C0 \sr_54_[12]  (.D(\sr_53_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[12]_net_1 ));
    DFN1E1C0 \sr_35_[5]  (.D(\sr_34_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[5]_net_1 ));
    DFN1E1C0 \sr_15_[12]  (.D(\sr_14_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[12]_net_1 ));
    DFN1E1C0 \sr_32_[6]  (.D(\sr_31_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[6]_net_1 ));
    DFN1E1C0 \sr_26_[12]  (.D(\sr_25_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[12]_net_1 ));
    DFN1E1C0 \sr_35_[4]  (.D(\sr_34_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[4]_net_1 ));
    DFN1E1C0 \sr_26_[9]  (.D(\sr_25_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[9]_net_1 ));
    DFN1E1C0 \sr_24_[12]  (.D(\sr_23_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[12]_net_1 ));
    DFN1E1C0 \sr_51_[4]  (.D(\sr_50_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[4]_net_1 ));
    DFN1E1C0 \sr_10_[7]  (.D(\sr_9_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[7]_net_1 ));
    DFN1E1C0 \sr_8_[2]  (.D(\sr_7_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[2]_net_1 ));
    DFN1E1C0 \sr_40_[12]  (.D(\sr_39_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[12]_net_1 ));
    DFN1E1C0 \sr_8_[8]  (.D(\sr_7_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[8]_net_1 ));
    DFN1E1C0 \sr_26_[1]  (.D(\sr_25_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[1]_net_1 ));
    DFN1E1C0 \sr_61_[4]  (.D(\sr_60_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[4]_net_1 ));
    DFN1E1C0 \sr_0_[0]  (.D(cur_error[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[0]));
    DFN1E1C0 \sr_43_[6]  (.D(\sr_42_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[6]_net_1 ));
    DFN1E1C0 \sr_10_[6]  (.D(\sr_9_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[6]_net_1 ));
    DFN1E1C0 \sr_21_[7]  (.D(\sr_20_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[7]_net_1 ));
    DFN1E1C0 \sr_0_[6]  (.D(cur_error[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[6]));
    DFN1E1C0 \sr_40_[5]  (.D(\sr_39_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[5]_net_1 ));
    DFN1E1C0 \sr_40_[10]  (.D(\sr_39_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[10]_net_1 ));
    DFN1E1C0 \sr_43_[10]  (.D(\sr_42_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[10]_net_1 ));
    DFN1E1C0 \sr_38_[1]  (.D(\sr_37_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[1]_net_1 ));
    DFN1E1C0 \sr_49_[1]  (.D(\sr_48_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[1]_net_1 ));
    DFN1E1C0 \sr_63_[11]  (.D(\sr_62_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[11]));
    DFN1E1C0 \sr_20_[9]  (.D(\sr_19_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[9]_net_1 ));
    DFN1E1C0 \sr_38_[2]  (.D(\sr_37_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[2]_net_1 ));
    DFN1E1C0 \sr_38_[7]  (.D(\sr_37_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[7]_net_1 ));
    DFN1E1C0 \sr_52_[1]  (.D(\sr_51_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[1]_net_1 ));
    DFN1E1C0 \sr_20_[1]  (.D(\sr_19_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[1]_net_1 ));
    DFN1E1C0 \sr_1_[0]  (.D(sr_new[0]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[0]));
    DFN1E1C0 \sr_61_[9]  (.D(\sr_60_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[9]_net_1 ));
    DFN1E1C0 \sr_0_[1]  (.D(cur_error[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[1]));
    DFN1E1C0 \sr_15_[4]  (.D(\sr_14_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[4]_net_1 ));
    DFN1E1C0 \sr_1_[6]  (.D(sr_new[6]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[6]));
    DFN1E1C0 \sr_62_[1]  (.D(\sr_61_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[1]_net_1 ));
    DFN1E1C0 \sr_25_[8]  (.D(\sr_24_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[8]_net_1 ));
    DFN1E1C0 \sr_48_[9]  (.D(\sr_47_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[9]_net_1 ));
    DFN1E1C0 \sr_1_[11]  (.D(sr_new[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_prev[11]));
    DFN1E1C0 \sr_49_[10]  (.D(\sr_48_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[10]_net_1 ));
    DFN1E1C0 \sr_53_[12]  (.D(\sr_52_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[12]_net_1 ));
    DFN1E1C0 \sr_13_[1]  (.D(\sr_12_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[1]_net_1 ));
    DFN1E1C0 \sr_7_[5]  (.D(\sr_6_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[5]_net_1 ));
    DFN1E1C0 \sr_5_[12]  (.D(\sr_4_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[12]_net_1 ));
    DFN1E1C0 \sr_47_[1]  (.D(\sr_46_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[1]_net_1 ));
    DFN1E1C0 \sr_23_[12]  (.D(\sr_22_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[12]_net_1 ));
    DFN1E1C0 \sr_63_[5]  (.D(\sr_62_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[5]));
    DFN1E1C0 \sr_45_[2]  (.D(\sr_44_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[2]_net_1 ));
    DFN1E1C0 \sr_2_[2]  (.D(sr_prev[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[2]_net_1 ));
    DFN1E1C0 \sr_2_[8]  (.D(sr_prev[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[8]_net_1 ));
    DFN1E1C0 \sr_11_[9]  (.D(\sr_10_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[9]_net_1 ));
    DFN1E1C0 \sr_33_[5]  (.D(\sr_32_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[5]_net_1 ));
    DFN1E1C0 \sr_59_[2]  (.D(\sr_58_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[2]_net_1 ));
    DFN1E1C0 \sr_12_[7]  (.D(\sr_11_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[7]_net_1 ));
    DFN1E1C0 \sr_6_[0]  (.D(\sr_5_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[0]_net_1 ));
    DFN1E1C0 \sr_41_[0]  (.D(\sr_40_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[0]_net_1 ));
    DFN1E1C0 \sr_1_[1]  (.D(sr_new[1]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[1]));
    DFN1E1C0 \sr_33_[4]  (.D(\sr_32_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[4]_net_1 ));
    DFN1E1C0 \sr_9_[12]  (.D(\sr_8_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[12]_net_1 ));
    DFN1E1C0 \sr_25_[0]  (.D(\sr_24_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[0]_net_1 ));
    DFN1E1C0 \sr_6_[6]  (.D(\sr_5_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[6]_net_1 ));
    DFN1E1C0 \sr_15_[10]  (.D(\sr_14_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[10]_net_1 ));
    DFN1E1C0 \sr_12_[6]  (.D(\sr_11_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[6]_net_1 ));
    DFN1E1C0 \sr_61_[3]  (.D(\sr_60_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[3]_net_1 ));
    DFN1E1C0 \sr_5_[0]  (.D(\sr_4_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[0]_net_1 ));
    DFN1E1C0 \sr_44_[3]  (.D(\sr_43_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[3]_net_1 ));
    DFN1E1C0 \sr_38_[0]  (.D(\sr_37_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[0]_net_1 ));
    DFN1E1C0 \sr_42_[5]  (.D(\sr_41_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[5]_net_1 ));
    DFN1E1C0 \sr_5_[6]  (.D(\sr_4_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[6]_net_1 ));
    DFN1E1C0 \sr_3_[5]  (.D(\sr_2_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[5]_net_1 ));
    DFN1E1C0 \sr_4_[3]  (.D(\sr_3_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[3]_net_1 ));
    DFN1E1C0 \sr_9_[9]  (.D(\sr_8_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[9]_net_1 ));
    DFN1E1C0 \sr_37_[10]  (.D(\sr_36_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[10]_net_1 ));
    DFN1E1C0 \sr_22_[9]  (.D(\sr_21_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[9]_net_1 ));
    DFN1E1C0 \sr_59_[4]  (.D(\sr_58_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[4]_net_1 ));
    DFN1E1C0 \sr_16_[10]  (.D(\sr_15_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[10]_net_1 ));
    DFN1E1C0 \sr_57_[2]  (.D(\sr_56_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[2]_net_1 ));
    DFN1E1C0 \sr_46_[3]  (.D(\sr_45_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[3]_net_1 ));
    DFN1E1C0 \sr_6_[1]  (.D(\sr_5_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[1]_net_1 ));
    DFN1E1C0 \sr_45_[8]  (.D(\sr_44_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[8]_net_1 ));
    DFN1E1C0 \sr_22_[1]  (.D(\sr_21_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[1]_net_1 ));
    DFN1E1C0 \sr_29_[7]  (.D(\sr_28_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[7]_net_1 ));
    DFN1E1C0 \sr_11_[12]  (.D(\sr_10_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[12]_net_1 ));
    DFN1E1C0 \sr_5_[1]  (.D(\sr_4_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[1]_net_1 ));
    DFN1E1C0 \sr_4_[10]  (.D(\sr_3_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[10]_net_1 ));
    DFN1E1C0 \sr_55_[3]  (.D(\sr_54_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[3]_net_1 ));
    DFN1E1C0 \sr_25_[2]  (.D(\sr_24_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[2]_net_1 ));
    DFN1E1C0 \sr_13_[4]  (.D(\sr_12_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[4]_net_1 ));
    DFN1E1C0 \sr_62_[10]  (.D(\sr_61_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[10]_net_1 ));
    DFN1E1C0 \sr_23_[8]  (.D(\sr_22_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[8]_net_1 ));
    DFN1E1C0 \sr_25_[5]  (.D(\sr_24_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[5]_net_1 ));
    DFN1E1C0 \sr_15_[8]  (.D(\sr_14_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[8]_net_1 ));
    DFN1E1C0 \sr_34_[10]  (.D(\sr_33_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[10]_net_1 ));
    DFN1E1C0 \sr_57_[4]  (.D(\sr_56_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[4]_net_1 ));
    DFN1E1C0 \sr_40_[3]  (.D(\sr_39_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[3]_net_1 ));
    DFN1E1C0 \sr_48_[4]  (.D(\sr_47_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[4]_net_1 ));
    DFN1E1C0 \sr_38_[3]  (.D(\sr_37_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[3]_net_1 ));
    DFN1E1C0 \sr_43_[2]  (.D(\sr_42_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[2]_net_1 ));
    DFN1E1C0 \sr_58_[6]  (.D(\sr_57_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[6]_net_1 ));
    DFN1E1C0 \sr_54_[9]  (.D(\sr_53_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[9]_net_1 ));
    DFN1E1C0 \sr_28_[4]  (.D(\sr_27_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[4]_net_1 ));
    DFN1E1C0 \sr_27_[7]  (.D(\sr_26_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[7]_net_1 ));
    DFN1E1C0 \sr_24_[6]  (.D(\sr_23_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[6]_net_1 ));
    DFN1E1C0 \sr_40_[11]  (.D(\sr_39_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[11]_net_1 ));
    DFN1E1C0 \sr_11_[10]  (.D(\sr_10_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[10]_net_1 ));
    DFN1E1C0 \sr_23_[0]  (.D(\sr_22_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[0]_net_1 ));
    DFN1E1C0 \sr_11_[11]  (.D(\sr_10_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[11]_net_1 ));
    DFN1E1C0 \sr_59_[12]  (.D(\sr_58_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[12]_net_1 ));
    DFN1E1C0 \sr_8_[9]  (.D(\sr_7_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[9]_net_1 ));
    DFN1E1C0 \sr_1_[10]  (.D(sr_new[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_prev[10]));
    DFN1E1C0 \sr_41_[7]  (.D(\sr_40_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[7]_net_1 ));
    DFN1E1C0 \sr_29_[12]  (.D(\sr_28_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[12]_net_1 ));
    DFN1E1C0 \sr_19_[9]  (.D(\sr_18_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[9]_net_1 ));
    DFN1E1C0 \sr_56_[9]  (.D(\sr_55_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[9]_net_1 ));
    DFN1E1C0 \sr_51_[7]  (.D(\sr_50_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[7]_net_1 ));
    DFN1E1C0 \sr_39_[11]  (.D(\sr_38_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[11]_net_1 ));
    DFN1E1C0 \sr_26_[6]  (.D(\sr_25_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[6]_net_1 ));
    DFN1E1C0 \sr_51_[8]  (.D(\sr_50_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[8]_net_1 ));
    DFN1E1C0 \sr_50_[12]  (.D(\sr_49_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[12]_net_1 ));
    DFN1E1C0 \sr_49_[0]  (.D(\sr_48_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[0]_net_1 ));
    DFN1E1C0 \sr_0_[5]  (.D(cur_error[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[5]));
    DFN1E1C0 \sr_15_[2]  (.D(\sr_14_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[2]_net_1 ));
    DFN1E1C0 \sr_61_[7]  (.D(\sr_60_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[7]_net_1 ));
    DFN1E1C0 \sr_48_[6]  (.D(\sr_47_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[6]_net_1 ));
    DFN1E1C0 \sr_15_[0]  (.D(\sr_14_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[0]_net_1 ));
    DFN1E1C0 \sr_35_[8]  (.D(\sr_34_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[8]_net_1 ));
    DFN1E1C0 \sr_61_[8]  (.D(\sr_60_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[8]_net_1 ));
    DFN1E1C0 \sr_20_[12]  (.D(\sr_19_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[12]_net_1 ));
    DFN1E1C0 \sr_43_[8]  (.D(\sr_42_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[8]_net_1 ));
    DFN1E1C0 \sr_11_[5]  (.D(\sr_10_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[5]_net_1 ));
    DFN1E1C0 \sr_50_[10]  (.D(\sr_49_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[10]_net_1 ));
    DFN1E1C0 \sr_55_[5]  (.D(\sr_54_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[5]_net_1 ));
    DFN1E1C0 \sr_53_[10]  (.D(\sr_52_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[10]_net_1 ));
    DFN1E1C0 \sr_48_[12]  (.D(\sr_47_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[12]_net_1 ));
    DFN1E1C0 \sr_32_[12]  (.D(\sr_31_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[12]_net_1 ));
    DFN1E1C0 \sr_11_[3]  (.D(\sr_10_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[3]_net_1 ));
    DFN1E1C0 \sr_0_[11]  (.D(cur_error[11]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable), .Q(sr_new[11]));
    DFN1E1C0 \sr_20_[10]  (.D(\sr_19_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[10]_net_1 ));
    DFN1E1C0 \sr_50_[9]  (.D(\sr_49_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[9]_net_1 ));
    DFN1E1C0 \sr_17_[9]  (.D(\sr_16_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[9]_net_1 ));
    DFN1E1C0 \sr_23_[10]  (.D(\sr_22_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[10]_net_1 ));
    DFN1E1C0 \sr_20_[6]  (.D(\sr_19_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[6]_net_1 ));
    DFN1E1C0 \sr_53_[3]  (.D(\sr_52_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[3]_net_1 ));
    DFN1E1C0 \sr_23_[2]  (.D(\sr_22_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[2]_net_1 ));
    DFN1E1C0 \sr_1_[5]  (.D(sr_new[5]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[5]));
    DFN1E1C0 \sr_61_[0]  (.D(\sr_60_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[0]_net_1 ));
    DFN1E1C0 \sr_47_[0]  (.D(\sr_46_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[0]_net_1 ));
    DFN1E1C0 \sr_23_[5]  (.D(\sr_22_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[5]_net_1 ));
    DFN1E1C0 \sr_42_[3]  (.D(\sr_41_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[3]_net_1 ));
    DFN1E1C0 \sr_25_[3]  (.D(\sr_24_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[3]_net_1 ));
    DFN1E1C0 \sr_35_[9]  (.D(\sr_34_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[9]_net_1 ));
    DFN1E1C0 \sr_13_[8]  (.D(\sr_12_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[8]_net_1 ));
    DFN1E1C0 \sr_36_[11]  (.D(\sr_35_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[11]_net_1 ));
    DFN1E1C0 \sr_51_[0]  (.D(\sr_50_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[0]_net_1 ));
    DFN1E1C0 \sr_18_[1]  (.D(\sr_17_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[1]_net_1 ));
    DFN1E1C0 \sr_2_[9]  (.D(sr_prev[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[9]_net_1 ));
    DFN1E1C0 \sr_9_[0]  (.D(\sr_8_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[0]_net_1 ));
    DFN1E1C0 \sr_59_[10]  (.D(\sr_58_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[10]_net_1 ));
    DFN1E1C0 \sr_35_[11]  (.D(\sr_34_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[11]_net_1 ));
    DFN1E1C0 \sr_35_[6]  (.D(\sr_34_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[6]_net_1 ));
    DFN1E1C0 \sr_9_[6]  (.D(\sr_8_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[6]_net_1 ));
    DFN1E1C0 \sr_29_[10]  (.D(\sr_28_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[10]_net_1 ));
    DFN1E1C0 \sr_44_[1]  (.D(\sr_43_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[1]_net_1 ));
    DFN1E1C0 \sr_38_[5]  (.D(\sr_37_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[5]_net_1 ));
    DFN1E1C0 \sr_37_[12]  (.D(\sr_36_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[12]_net_1 ));
    DFN1E1C0 \sr_6_[5]  (.D(\sr_5_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[5]_net_1 ));
    DFN1E1C0 \sr_48_[11]  (.D(\sr_47_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[11]_net_1 ));
    DFN1E1C0 \sr_38_[4]  (.D(\sr_37_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[4]_net_1 ));
    DFN1E1C0 \sr_4_[4]  (.D(\sr_3_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[4]_net_1 ));
    DFN1E1C0 \sr_38_[10]  (.D(\sr_37_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[10]_net_1 ));
    DFN1E1C0 \sr_5_[5]  (.D(\sr_4_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[5]_net_1 ));
    DFN1E1C0 \sr_13_[2]  (.D(\sr_12_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[2]_net_1 ));
    DFN1E1C0 \sr_46_[1]  (.D(\sr_45_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[1]_net_1 ));
    DFN1E1C0 \sr_9_[1]  (.D(\sr_8_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[1]_net_1 ));
    DFN1E1C0 \sr_13_[0]  (.D(\sr_12_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[0]_net_1 ));
    DFN1E1C0 \sr_33_[8]  (.D(\sr_32_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[8]_net_1 ));
    DFN1E1C0 \sr_49_[7]  (.D(\sr_48_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[7]_net_1 ));
    DFN1E1C0 \sr_59_[7]  (.D(\sr_58_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[7]_net_1 ));
    DFN1E1C0 \sr_52_[9]  (.D(\sr_51_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[9]_net_1 ));
    DFN1E1C0 \sr_59_[8]  (.D(\sr_58_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[8]_net_1 ));
    DFN1E1C0 \sr_53_[5]  (.D(\sr_52_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[5]_net_1 ));
    DFN1E1C0 \sr_22_[6]  (.D(\sr_21_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[6]_net_1 ));
    DFN1E1C0 \sr_55_[1]  (.D(\sr_54_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[1]_net_1 ));
    DFN1E1C0 \sr_54_[2]  (.D(\sr_53_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[2]_net_1 ));
    DFN1E1C0 \sr_43_[11]  (.D(\sr_42_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[11]_net_1 ));
    DFN1E1C0 \sr_8_[0]  (.D(\sr_7_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[0]_net_1 ));
    DFN1E1C0 \sr_23_[3]  (.D(\sr_22_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[3]_net_1 ));
    DFN1E1C0 \sr_40_[1]  (.D(\sr_39_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[1]_net_1 ));
    DFN1E1C0 \sr_33_[9]  (.D(\sr_32_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[9]_net_1 ));
    DFN1E1C0 \sr_19_[5]  (.D(\sr_18_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[5]_net_1 ));
    DFN1E1C0 \sr_18_[4]  (.D(\sr_17_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[4]_net_1 ));
    DFN1E1C0 \sr_28_[8]  (.D(\sr_27_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[8]_net_1 ));
    DFN1E1C0 \sr_8_[6]  (.D(\sr_7_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[6]_net_1 ));
    DFN1E1C0 \sr_32_[11]  (.D(\sr_31_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[11]_net_1 ));
    DFN1E1C0 \sr_61_[12]  (.D(\sr_60_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[12]_net_1 ));
    DFN1E1C0 \sr_19_[3]  (.D(\sr_18_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[3]_net_1 ));
    DFN1E1C0 \sr_8_[11]  (.D(\sr_7_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[11]_net_1 ));
    DFN1E1C0 \sr_47_[7]  (.D(\sr_46_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[7]_net_1 ));
    DFN1E1C0 \sr_57_[7]  (.D(\sr_56_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[7]_net_1 ));
    DFN1E1C0 \sr_56_[2]  (.D(\sr_55_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[2]_net_1 ));
    DFN1E1C0 \sr_17_[10]  (.D(\sr_16_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[10]_net_1 ));
    DFN1E1C0 \sr_57_[8]  (.D(\sr_56_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[8]_net_1 ));
    DFN1E1C0 \sr_48_[2]  (.D(\sr_47_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[2]_net_1 ));
    DFN1E1C0 \sr_15_[7]  (.D(\sr_14_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[7]_net_1 ));
    DFN1E1C0 \sr_34_[11]  (.D(\sr_33_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[11]_net_1 ));
    DFN1E1C0 \sr_33_[6]  (.D(\sr_32_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[6]_net_1 ));
    DFN1E1C0 \sr_54_[4]  (.D(\sr_53_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[4]_net_1 ));
    DFN1E1C0 \sr_15_[6]  (.D(\sr_14_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[6]_net_1 ));
    DFN1E1C0 \sr_59_[0]  (.D(\sr_58_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[0]_net_1 ));
    DFN1E1C0 \sr_50_[11]  (.D(\sr_49_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[11]_net_1 ));
    DFN1E1C0 \sr_45_[5]  (.D(\sr_44_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[5]_net_1 ));
    DFN1E1C0 \sr_8_[1]  (.D(\sr_7_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[1]_net_1 ));
    DFN1E1C0 \sr_31_[1]  (.D(\sr_30_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[1]_net_1 ));
    DFN1E1C0 \sr_28_[0]  (.D(\sr_27_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[0]_net_1 ));
    DFN1E1C0 \sr_17_[5]  (.D(\sr_16_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[5]_net_1 ));
    DFN1E1C0 \sr_24_[7]  (.D(\sr_23_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[7]_net_1 ));
    DFN1E1C0 \sr_20_[11]  (.D(\sr_19_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[11]_net_1 ));
    DFN1E1C0 \sr_31_[2]  (.D(\sr_30_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[2]_net_1 ));
    DFN1E1C0 \sr_17_[3]  (.D(\sr_16_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[3]_net_1 ));
    DFN1E1C0 \sr_56_[4]  (.D(\sr_55_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[4]_net_1 ));
    DFN1E1C0 \sr_31_[7]  (.D(\sr_30_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[7]_net_1 ));
    DFN1E1C0 \sr_25_[9]  (.D(\sr_24_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[9]_net_1 ));
    DFN1E1C0 \sr_61_[10]  (.D(\sr_60_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[10]_net_1 ));
    DFN1E1C0 \sr_50_[2]  (.D(\sr_49_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[2]_net_1 ));
    DFN1E1C0 \sr_14_[10]  (.D(\sr_13_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[10]_net_1 ));
    DFN1E1C0 \sr_61_[11]  (.D(\sr_60_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[11]_net_1 ));
    DFN1E1C0 \sr_25_[1]  (.D(\sr_24_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[1]_net_1 ));
    DFN1E1C0 \sr_60_[2]  (.D(\sr_59_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[2]_net_1 ));
    DFN1E1C0 \sr_26_[7]  (.D(\sr_25_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[7]_net_1 ));
    DFN1E1C0 \sr_2_[0]  (.D(sr_prev[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[0]_net_1 ));
    DFN1E1C0 \sr_41_[9]  (.D(\sr_40_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[9]_net_1 ));
    DFN1E1C0 \sr_57_[0]  (.D(\sr_56_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[0]_net_1 ));
    DFN1E1C0 \sr_48_[8]  (.D(\sr_47_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[8]_net_1 ));
    DFN1E1C0 \sr_53_[1]  (.D(\sr_52_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[1]_net_1 ));
    DFN1E1C0 \sr_2_[6]  (.D(sr_prev[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[6]_net_1 ));
    DFN1E1C0 \sr_7_[7]  (.D(\sr_6_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[7]_net_1 ));
    DFN1E1C0 \sr_42_[1]  (.D(\sr_41_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[1]_net_1 ));
    DFN1E1C0 \sr_63_[1]  (.D(\sr_62_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[1]));
    DFN1E1C0 \sr_50_[4]  (.D(\sr_49_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[4]_net_1 ));
    DFN1E1C0 \sr_58_[12]  (.D(\sr_57_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[12]_net_1 ));
    DFN1E1C0 \sr_58_[3]  (.D(\sr_57_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[3]_net_1 ));
    DFN1E1C0 \sr_28_[2]  (.D(\sr_27_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[2]_net_1 ));
    DFN1E1C0 \sr_4_[2]  (.D(\sr_3_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[2]_net_1 ));
    DFN1E1C0 \sr_4_[8]  (.D(\sr_3_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[8]_net_1 ));
    DFN1E1C0 \sr_28_[5]  (.D(\sr_27_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[5]_net_1 ));
    DFN1E1C0 \sr_28_[12]  (.D(\sr_27_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[12]_net_1 ));
    DFN1E1C0 \sr_60_[4]  (.D(\sr_59_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[4]_net_1 ));
    DFN1E1C0 \sr_19_[11]  (.D(\sr_18_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[11]_net_1 ));
    DFN1E1C0 \sr_14_[9]  (.D(\sr_13_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[9]_net_1 ));
    DFN1E1C0 \sr_18_[8]  (.D(\sr_17_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[8]_net_1 ));
    DFN1E1C0 \sr_47_[11]  (.D(\sr_46_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[11]_net_1 ));
    DFN1E1C0 \sr_20_[7]  (.D(\sr_19_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[7]_net_1 ));
    DFN1E1C0 \sr_2_[1]  (.D(sr_prev[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[1]_net_1 ));
    DFN1E1C0 \sr_31_[0]  (.D(\sr_30_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[0]_net_1 ));
    DFN1E1C0 \sr_42_[10]  (.D(\sr_41_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[10]_net_1 ));
    DFN1E1C0 \sr_44_[0]  (.D(\sr_43_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[0]_net_1 ));
    DFN1E1C0 \sr_13_[7]  (.D(\sr_12_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[7]_net_1 ));
    DFN1E1C0 \sr_36_[12]  (.D(\sr_35_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[12]_net_1 ));
    DFN1E1C0 \sr_9_[5]  (.D(\sr_8_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[5]_net_1 ));
    DFN1E1C0 \sr_34_[12]  (.D(\sr_33_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[12]_net_1 ));
    DFN1E1C0 \sr_3_[7]  (.D(\sr_2_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[7]_net_1 ));
    DFN1E1C0 \sr_13_[6]  (.D(\sr_12_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[6]_net_1 ));
    DFN1E1C0 \sr_16_[9]  (.D(\sr_15_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[9]_net_1 ));
    DFN1E1C0 \sr_12_[12]  (.D(\sr_11_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[12]_net_1 ));
    DFN1E1C0 \sr_43_[5]  (.D(\sr_42_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[5]_net_1 ));
    DFN1E1C0 \sr_46_[0]  (.D(\sr_45_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[0]_net_1 ));
    DFN1E1C0 \sr_52_[2]  (.D(\sr_51_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[2]_net_1 ));
    DFN1E1C0 \sr_60_[9]  (.D(\sr_59_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[9]_net_1 ));
    DFN1E1C0 \sr_4_[12]  (.D(\sr_3_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[12]_net_1 ));
    DFN1E1C0 \sr_58_[11]  (.D(\sr_57_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[11]_net_1 ));
    DFN1E1C0 \sr_3_[12]  (.D(\sr_2_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[12]_net_1 ));
    DFN1E1C0 \sr_23_[9]  (.D(\sr_22_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[9]_net_1 ));
    DFN1E1C0 \sr_28_[11]  (.D(\sr_27_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[11]_net_1 ));
    DFN1E1C0 \sr_62_[2]  (.D(\sr_61_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[2]_net_1 ));
    DFN1E1C0 \sr_16_[11]  (.D(\sr_15_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[11]_net_1 ));
    DFN1E1C0 \sr_1_[12]  (.D(sr_new_0_0), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_prev[12]));
    DFN1E1C0 \sr_18_[2]  (.D(\sr_17_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[2]_net_1 ));
    DFN1E1C0 \sr_39_[1]  (.D(\sr_38_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[1]_net_1 ));
    DFN1E1C0 \sr_23_[1]  (.D(\sr_22_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[1]_net_1 ));
    DFN1E1C0 \sr_18_[0]  (.D(\sr_17_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[0]_net_1 ));
    DFN1E1C0 \sr_38_[8]  (.D(\sr_37_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[8]_net_1 ));
    DFN1E1C0 \sr_8_[10]  (.D(\sr_7_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[10]_net_1 ));
    DFN1E1C0 \sr_10_[9]  (.D(\sr_9_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[9]_net_1 ));
    DFN1E1C0 \sr_45_[12]  (.D(\sr_44_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[12]_net_1 ));
    DFN1E1C0 \sr_39_[2]  (.D(\sr_38_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[2]_net_1 ));
    DFN1E1C0 \sr_8_[12]  (.D(\sr_7_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[12]_net_1 ));
    DFN1E1C0 \sr_15_[11]  (.D(\sr_14_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[11]_net_1 ));
    DFN1E1C0 \sr_39_[7]  (.D(\sr_38_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[7]_net_1 ));
    DFN1E1C0 \sr_52_[4]  (.D(\sr_51_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[4]_net_1 ));
    DFN1E1C0 \sr_41_[4]  (.D(\sr_40_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[4]_net_1 ));
    DFN1E1C0 \sr_58_[5]  (.D(\sr_57_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[5]_net_1 ));
    DFN1E1C0 \sr_40_[0]  (.D(\sr_39_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[0]_net_1 ));
    DFN1E1C0 \sr_31_[3]  (.D(\sr_30_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[3]_net_1 ));
    DFN1E1C0 \sr_51_[6]  (.D(\sr_50_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[6]_net_1 ));
    DFN1E1C0 \sr_17_[12]  (.D(\sr_16_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[12]_net_1 ));
    DFN1E1C0 \sr_45_[3]  (.D(\sr_44_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[3]_net_1 ));
    DFN1E1C0 \sr_62_[4]  (.D(\sr_61_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[4]_net_1 ));
    DFN1E1C0 \sr_21_[4]  (.D(\sr_20_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[4]_net_1 ));
    DFN1E1C0 \sr_60_[3]  (.D(\sr_59_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[3]_net_1 ));
    DFN1E1C0 \sr_22_[7]  (.D(\sr_21_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[7]_net_1 ));
    DFN1E1C0 \sr_61_[6]  (.D(\sr_60_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[6]_net_1 ));
    DFN1E1C0 \sr_49_[9]  (.D(\sr_48_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[9]_net_1 ));
    DFN1E1C0 \sr_18_[10]  (.D(\sr_17_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[10]_net_1 ));
    DFN1E1C0 \sr_8_[5]  (.D(\sr_7_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[5]_net_1 ));
    DFN1E1C0 \sr_33_[12]  (.D(\sr_32_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[12]_net_1 ));
    DFN1E1C0 \sr_28_[3]  (.D(\sr_27_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[3]_net_1 ));
    DFN1E1C0 \sr_38_[9]  (.D(\sr_37_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[9]_net_1 ));
    DFN1E1C0 \sr_53_[11]  (.D(\sr_52_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[11]_net_1 ));
    DFN1E1C0 \sr_37_[1]  (.D(\sr_36_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[1]_net_1 ));
    DFN1E1C0 \sr_37_[2]  (.D(\sr_36_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[2]_net_1 ));
    DFN1E1C0 \sr_23_[11]  (.D(\sr_22_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[11]_net_1 ));
    DFN1E1C0 \sr_3_[11]  (.D(\sr_2_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[11]_net_1 ));
    DFN1E1C0 \sr_37_[7]  (.D(\sr_36_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[7]_net_1 ));
    DFN1E1C0 \sr_38_[6]  (.D(\sr_37_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[6]_net_1 ));
    DFN1E1C0 \sr_41_[6]  (.D(\sr_40_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[6]_net_1 ));
    DFN1E1C0 \sr_44_[7]  (.D(\sr_43_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[7]_net_1 ));
    DFN1E1C0 \sr_54_[7]  (.D(\sr_53_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[7]_net_1 ));
    DFN1E1C0 \sr_0_[7]  (.D(cur_error[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[7]));
    DFN1E1C0 \sr_9_[11]  (.D(\sr_8_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[11]_net_1 ));
    DFN1E1C0 \sr_62_[9]  (.D(\sr_61_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[9]_net_1 ));
    DFN1E1C0 \sr_54_[8]  (.D(\sr_53_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[8]_net_1 ));
    DFN1E1C0 \sr_39_[0]  (.D(\sr_38_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[0]_net_1 ));
    DFN1E1C0 \sr_47_[9]  (.D(\sr_46_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[9]_net_1 ));
    DFN1E1C0 \sr_6_[12]  (.D(\sr_5_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[12]_net_1 ));
    DFN1E1C0 \sr_7_[11]  (.D(\sr_6_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[11]_net_1 ));
    DFN1E1C0 \sr_46_[7]  (.D(\sr_45_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[7]_net_1 ));
    DFN1E1C0 \sr_14_[5]  (.D(\sr_13_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[5]_net_1 ));
    DFN1E1C0 \sr_56_[7]  (.D(\sr_55_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[7]_net_1 ));
    DFN1E1C0 \sr_12_[9]  (.D(\sr_11_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[9]_net_1 ));
    DFN1E1C0 \sr_12_[11]  (.D(\sr_11_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[11]_net_1 ));
    DFN1E1C0 \sr_55_[9]  (.D(\sr_54_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[9]_net_1 ));
    DFN1E1C0 \sr_56_[8]  (.D(\sr_55_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[8]_net_1 ));
    DFN1E1C0 \sr_25_[6]  (.D(\sr_24_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[6]_net_1 ));
    DFN1E1C0 \sr_14_[3]  (.D(\sr_13_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[3]_net_1 ));
    DFN1E1C0 \sr_42_[0]  (.D(\sr_41_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[0]_net_1 ));
    DFN1E1C0 \sr_1_[7]  (.D(sr_new[7]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[7]));
    DFN1E1C0 \sr_2_[5]  (.D(sr_prev[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[5]_net_1 ));
    DFN1E1C0 \sr_14_[11]  (.D(\sr_13_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[11]_net_1 ));
    DFN1E1C0 \sr_37_[0]  (.D(\sr_36_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[0]_net_1 ));
    DFN1E1C0 \sr_58_[1]  (.D(\sr_57_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[1]_net_1 ));
    DFN1E1C0 \sr_11_[1]  (.D(\sr_10_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[1]_net_1 ));
    DFN1E1C0 \sr_62_[3]  (.D(\sr_61_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[3]_net_1 ));
    DFN1E1C0 \sr_45_[10]  (.D(\sr_44_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[10]_net_1 ));
    DFN1E1C0 \sr_16_[5]  (.D(\sr_15_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[5]_net_1 ));
    DFN1E1C0 \sr_43_[3]  (.D(\sr_42_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[3]_net_1 ));
    DFN1E1C0 \sr_61_[5]  (.D(\sr_60_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[5]_net_1 ));
    DFN1E1C0 \sr_54_[0]  (.D(\sr_53_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[0]_net_1 ));
    DFN1E1C0 \sr_16_[3]  (.D(\sr_15_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[3]_net_1 ));
    DFN1E1C0 \sr_4_[9]  (.D(\sr_3_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[9]_net_1 ));
    DFN1E1C0 \sr_40_[7]  (.D(\sr_39_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[7]_net_1 ));
    DFN1E1C0 \sr_50_[7]  (.D(\sr_49_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[7]_net_1 ));
    DFN1E1C0 \sr_31_[5]  (.D(\sr_30_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[5]_net_1 ));
    DFN1E1C0 \sr_50_[8]  (.D(\sr_49_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[8]_net_1 ));
    DFN1E1C0 \sr_49_[4]  (.D(\sr_48_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[4]_net_1 ));
    DFN1E1C0 \sr_31_[4]  (.D(\sr_30_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[4]_net_1 ));
    DFN1E1C0 \sr_0_[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable), .Q(sr_new[12]));
    DFN1E1C0 \sr_39_[3]  (.D(\sr_38_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[3]_net_1 ));
    DFN1E1C0 \sr_6_[7]  (.D(\sr_5_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[7]_net_1 ));
    DFN1E1C0 \sr_60_[7]  (.D(\sr_59_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[7]_net_1 ));
    DFN1E1C0 \sr_59_[6]  (.D(\sr_58_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[6]_net_1 ));
    DFN1E1C0 \sr_7_[3]  (.D(\sr_6_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[3]_net_1 ));
    DFN1E1C0 \sr_46_[10]  (.D(\sr_45_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[10]_net_1 ));
    DFN1E1C0 \sr_60_[8]  (.D(\sr_59_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[8]_net_1 ));
    DFN1E1C0 \sr_29_[4]  (.D(\sr_28_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[4]_net_1 ));
    DFN1E1C0 \sr_57_[11]  (.D(\sr_56_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[11]_net_1 ));
    DFN1E1C0 \sr_56_[0]  (.D(\sr_55_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[0]_net_1 ));
    DFN1E1C0 \sr_5_[7]  (.D(\sr_4_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[7]_net_1 ));
    DFN1E1C0 \sr_18_[7]  (.D(\sr_17_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[7]_net_1 ));
    DFN1E1C0 \sr_10_[5]  (.D(\sr_9_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[5]_net_1 ));
    DFN1E1C0 \sr_41_[12]  (.D(\sr_40_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[12]_net_1 ));
    DFN1E1C0 \sr_52_[10]  (.D(\sr_51_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[10]_net_1 ));
    DFN1E1C0 \sr_27_[11]  (.D(\sr_26_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[11]_net_1 ));
    DFN1E1C0 \sr_39_[12]  (.D(\sr_38_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[12]_net_1 ));
    DFN1E1C0 \sr_18_[6]  (.D(\sr_17_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[6]_net_1 ));
    DFN1E1C0 \sr_22_[10]  (.D(\sr_21_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[10]_net_1 ));
    DFN1E1C0 \sr_10_[3]  (.D(\sr_9_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[3]_net_1 ));
    DFN1E1C0 \sr_48_[5]  (.D(\sr_47_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[5]_net_1 ));
    DFN1E1C0 \sr_60_[0]  (.D(\sr_59_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[0]_net_1 ));
    DFN1E1C0 \sr_47_[4]  (.D(\sr_46_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[4]_net_1 ));
    DFN1E1C0 \sr_30_[12]  (.D(\sr_29_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[12]_net_1 ));
    DFN1E1C0 \sr_37_[3]  (.D(\sr_36_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[3]_net_1 ));
    DFN1E1C0 \sr_57_[6]  (.D(\sr_56_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[6]_net_1 ));
    DFN1E1C0 \sr_49_[6]  (.D(\sr_48_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[6]_net_1 ));
    DFN1E1C0 \sr_3_[3]  (.D(\sr_2_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[3]_net_1 ));
    DFN1E1C0 \sr_28_[9]  (.D(\sr_27_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[9]_net_1 ));
    DFN1E1C0 \sr_27_[4]  (.D(\sr_26_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[4]_net_1 ));
    DFN1E1C0 \sr_62_[12]  (.D(\sr_61_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[12]_net_1 ));
    DFN1E1C0 \sr_50_[0]  (.D(\sr_49_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[0]_net_1 ));
    DFN1E1C0 \sr_53_[9]  (.D(\sr_52_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[9]_net_1 ));
    DFN1E1C0 \sr_23_[6]  (.D(\sr_22_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[6]_net_1 ));
    DFN1E1C0 \sr_28_[1]  (.D(\sr_27_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[1]_net_1 ));
    DFN1E1C0 \sr_11_[4]  (.D(\sr_10_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[4]_net_1 ));
    DFN1E1C0 \sr_30_[10]  (.D(\sr_29_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[10]_net_1 ));
    DFN1E1C0 \sr_21_[8]  (.D(\sr_20_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[8]_net_1 ));
    DFN1E1C0 \sr_16_[12]  (.D(\sr_15_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[12]_net_1 ));
    DFN1E1C0 \sr_41_[10]  (.D(\sr_40_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[10]_net_1 ));
    DFN1E1C0 \sr_45_[1]  (.D(\sr_44_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[1]_net_1 ));
    DFN1E1C0 \sr_33_[10]  (.D(\sr_32_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[10]_net_1 ));
    DFN1E1C0 \sr_14_[12]  (.D(\sr_13_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[12]_net_1 ));
    DFN1E1C0 \sr_41_[11]  (.D(\sr_40_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[11]_net_1 ));
    DFN1E1C0 \sr_55_[12]  (.D(\sr_54_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[12]_net_1 ));
    DFN1E1C0 \sr_42_[7]  (.D(\sr_41_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[7]_net_1 ));
    DFN1E1C0 \sr_52_[7]  (.D(\sr_51_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[7]_net_1 ));
    DFN1E1C0 \sr_41_[2]  (.D(\sr_40_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[2]_net_1 ));
    DFN1E1C0 \sr_52_[8]  (.D(\sr_51_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[8]_net_1 ));
    DFN1E1C0 \sr_25_[12]  (.D(\sr_24_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[12]_net_1 ));
    DFN1E1C0 \sr_47_[6]  (.D(\sr_46_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[6]_net_1 ));
    DFN1E1C0 \sr_62_[7]  (.D(\sr_61_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[7]_net_1 ));
    DFN1E1C0 \sr_62_[8]  (.D(\sr_61_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[8]_net_1 ));
    DFN1E1C0 \sr_19_[1]  (.D(\sr_18_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[1]_net_1 ));
    DFN1E1C0 \sr_21_[0]  (.D(\sr_20_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[0]_net_1 ));
    DFN1E1C0 \sr_39_[10]  (.D(\sr_38_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[10]_net_1 ));
    DFN1E1C0 \sr_12_[5]  (.D(\sr_11_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[5]_net_1 ));
    DFN1E1C0 \sr_0_[10]  (.D(cur_error[10]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable), .Q(sr_new[10]));
    DFN1E1C0 \sr_12_[3]  (.D(\sr_11_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[3]_net_1 ));
    DFN1E1C0 \sr_34_[1]  (.D(\sr_33_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[1]_net_1 ));
    DFN1E1C0 \sr_39_[5]  (.D(\sr_38_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[5]_net_1 ));
    DFN1E1C0 \sr_5_[11]  (.D(\sr_4_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[11]_net_1 ));
    DFN1E1C0 \sr_34_[2]  (.D(\sr_33_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[2]_net_1 ));
    DFN1E1C0 \sr_39_[4]  (.D(\sr_38_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[4]_net_1 ));
    DFN1E1C0 \sr_55_[2]  (.D(\sr_54_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[2]_net_1 ));
    DFN1E1C0 \sr_62_[0]  (.D(\sr_61_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[0]_net_1 ));
    DFN1E1C0 \sr_34_[7]  (.D(\sr_33_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[7]_net_1 ));
    DFN1E1C0 \sr_41_[8]  (.D(\sr_40_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[8]_net_1 ));
    DFN1E1C0 \sr_52_[0]  (.D(\sr_51_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[0]_net_1 ));
    DFN1E1C0 \sr_17_[1]  (.D(\sr_16_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[1]_net_1 ));
    DFN1E1C0 \sr_4_[0]  (.D(\sr_3_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[0]_net_1 ));
    DFN1E1C0 \sr_36_[1]  (.D(\sr_35_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[1]_net_1 ));
    DFN1E1C0 \sr_13_[12]  (.D(\sr_12_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[12]_net_1 ));
    DFN1E1C0 \sr_4_[6]  (.D(\sr_3_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[6]_net_1 ));
    DFN1E1C0 \sr_44_[9]  (.D(\sr_43_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[9]_net_1 ));
    DFN1E1C0 \sr_0_[3]  (.D(cur_error[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[3]));
    DFN1E1C0 \sr_36_[2]  (.D(\sr_35_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[2]_net_1 ));
    DFN1E1C0 \sr_51_[3]  (.D(\sr_50_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[3]_net_1 ));
    DFN1E1C0 \sr_36_[7]  (.D(\sr_35_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[7]_net_1 ));
    DFN1E1C0 \sr_21_[2]  (.D(\sr_20_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[2]_net_1 ));
    DFN1E1C0 \sr_37_[5]  (.D(\sr_36_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[5]_net_1 ));
    DFN1E1C0 \sr_55_[4]  (.D(\sr_54_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[4]_net_1 ));
    DFN1E1C0 \sr_21_[5]  (.D(\sr_20_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[5]_net_1 ));
    DFN1E1C0 \sr_43_[1]  (.D(\sr_42_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[1]_net_1 ));
    DFN1E1C0 \sr_11_[8]  (.D(\sr_10_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[8]_net_1 ));
    DFN1E1C0 \sr_37_[4]  (.D(\sr_36_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[4]_net_1 ));
    DFN1E1C0 \sr_62_[11]  (.D(\sr_61_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[11]_net_1 ));
    DFN1E1C0 \sr_46_[9]  (.D(\sr_45_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[9]_net_1 ));
    DFN1E1C0 \sr_25_[7]  (.D(\sr_24_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[7]_net_1 ));
    DFN1E1C0 \sr_48_[3]  (.D(\sr_47_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[3]_net_1 ));
    DFN1E1C0 \sr_30_[1]  (.D(\sr_29_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[1]_net_1 ));
    DFN1E1C0 \sr_4_[1]  (.D(\sr_3_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[1]_net_1 ));
    DFN1E1C0 \sr_55_[10]  (.D(\sr_54_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[10]_net_1 ));
    DFN1E1C0 \sr_19_[4]  (.D(\sr_18_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[4]_net_1 ));
    DFN1E1C0 \sr_9_[7]  (.D(\sr_8_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[7]_net_1 ));
    DFN1E1C0 \sr_7_[4]  (.D(\sr_6_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[4]_net_1 ));
    DFN1E1C0 \sr_29_[8]  (.D(\sr_28_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[8]_net_1 ));
    DFN1E1C0 \sr_1_[3]  (.D(sr_new[3]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[3]));
    DFN1E1C0 \sr_34_[0]  (.D(\sr_33_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[0]_net_1 ));
    DFN1E1C0 \sr_30_[2]  (.D(\sr_29_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[2]_net_1 ));
    DFN1E1C0 \sr_25_[10]  (.D(\sr_24_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[10]_net_1 ));
    DFN1E1C0 \sr_30_[7]  (.D(\sr_29_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[7]_net_1 ));
    DFN1E1C0 \sr_49_[2]  (.D(\sr_48_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[2]_net_1 ));
    DFN1E1C0 \sr_56_[10]  (.D(\sr_55_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[10]_net_1 ));
    DFN1E1C0 \sr_40_[9]  (.D(\sr_39_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[9]_net_1 ));
    DFN1E1C0 \sr_36_[0]  (.D(\sr_35_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[0]_net_1 ));
    DFN1E1C0 \sr_11_[2]  (.D(\sr_10_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[2]_net_1 ));
    DFN1E1C0 \sr_30_[11]  (.D(\sr_29_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[11]_net_1 ));
    DFN1E1C0 \sr_53_[2]  (.D(\sr_52_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[2]_net_1 ));
    DFN1E1C0 \sr_26_[10]  (.D(\sr_25_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[10]_net_1 ));
    DFN1E1C0 \sr_11_[0]  (.D(\sr_10_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[0]_net_1 ));
    DFN1E1C0 \sr_31_[8]  (.D(\sr_30_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[8]_net_1 ));
    DFN1E1C0 \sr_29_[0]  (.D(\sr_28_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[0]_net_1 ));
    DFN1E1C0 \sr_17_[4]  (.D(\sr_16_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[4]_net_1 ));
    DFN1E1C0 \sr_6_[3]  (.D(\sr_5_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[3]_net_1 ));
    DFN1E1C0 \sr_51_[12]  (.D(\sr_50_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[12]_net_1 ));
    DFN1E1C0 \sr_27_[8]  (.D(\sr_26_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[8]_net_1 ));
    DFN1E1C0 \sr_3_[4]  (.D(\sr_2_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[4]_net_1 ));
    DFN1E1C0 \sr_63_[2]  (.D(\sr_62_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[2]));
    DFN1E1C0 \sr_21_[12]  (.D(\sr_20_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[12]_net_1 ));
    DFN1E1C0 \sr_5_[3]  (.D(\sr_4_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[3]_net_1 ));
    DFN1E1C0 \sr_15_[9]  (.D(\sr_14_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[9]_net_1 ));
    DFN1E1C0 \sr_51_[5]  (.D(\sr_50_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[5]_net_1 ));
    DFN1E1C0 \sr_47_[2]  (.D(\sr_46_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[2]_net_1 ));
    DFN1E1C0 \sr_47_[10]  (.D(\sr_46_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[10]_net_1 ));
    DFN1E1C0 \sr_45_[0]  (.D(\sr_44_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[0]_net_1 ));
    DFN1E1C0 \sr_58_[9]  (.D(\sr_57_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[9]_net_1 ));
    DFN1E1C0 \sr_30_[0]  (.D(\sr_29_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[0]_net_1 ));
    DFN1E1C0 \sr_44_[4]  (.D(\sr_43_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[4]_net_1 ));
    DFN1E1C0 \sr_53_[4]  (.D(\sr_52_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[4]_net_1 ));
    DFN1E1C0 \sr_34_[3]  (.D(\sr_33_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[3]_net_1 ));
    DFN1E1C0 \sr_54_[6]  (.D(\sr_53_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[6]_net_1 ));
    DFN1E1C0 \sr_49_[8]  (.D(\sr_48_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[8]_net_1 ));
    DFN1E1C0 \sr_28_[6]  (.D(\sr_27_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[6]_net_1 ));
    DFN1E1C0 \sr_21_[3]  (.D(\sr_20_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[3]_net_1 ));
    DFN1E1C0 \sr_31_[9]  (.D(\sr_30_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[9]_net_1 ));
    DFN1E1C0 \sr_8_[7]  (.D(\sr_7_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[7]_net_1 ));
    DFN1E1C0 \sr_27_[0]  (.D(\sr_26_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[0]_net_1 ));
    DFN1E1C0 \sr_24_[4]  (.D(\sr_23_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[4]_net_1 ));
    DFN1E1C0 \sr_63_[4]  (.D(\sr_62_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[4]));
    DFN1E1C0 \sr_32_[1]  (.D(\sr_31_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[1]_net_1 ));
    DFN1E1C0 \sr_19_[12]  (.D(\sr_18_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[12]_net_1 ));
    DFN1E1C0 \sr_23_[7]  (.D(\sr_22_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[7]_net_1 ));
    DFN1E1C0 \sr_51_[10]  (.D(\sr_50_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[10]_net_1 ));
    DFN1E1C0 \sr_32_[2]  (.D(\sr_31_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[2]_net_1 ));
    DFN1E1C0 \sr_38_[12]  (.D(\sr_37_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[12]_net_1 ));
    DFN1E1C0 \sr_59_[3]  (.D(\sr_58_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[3]_net_1 ));
    DFN1E1C0 \sr_51_[11]  (.D(\sr_50_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[11]_net_1 ));
    DFN1E1C0 \sr_29_[2]  (.D(\sr_28_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[2]_net_1 ));
    DFN1E1C0 \sr_32_[7]  (.D(\sr_31_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[7]_net_1 ));
    DFN1E1C0 \sr_21_[10]  (.D(\sr_20_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[10]_net_1 ));
    DFN1E1C0 \sr_46_[4]  (.D(\sr_45_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[4]_net_1 ));
    DFN1E1C0 \sr_31_[6]  (.D(\sr_30_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[6]_net_1 ));
    DFN1E1C0 \sr_36_[3]  (.D(\sr_35_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[3]_net_1 ));
    DFN1E1C0 \sr_29_[5]  (.D(\sr_28_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[5]_net_1 ));
    DFN1E1C0 \sr_56_[6]  (.D(\sr_55_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[6]_net_1 ));
    DFN1E1C0 \sr_21_[11]  (.D(\sr_20_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[11]_net_1 ));
    DFN1E1C0 \sr_19_[8]  (.D(\sr_18_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[8]_net_1 ));
    DFN1E1C0 \sr_44_[10]  (.D(\sr_43_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[10]_net_1 ));
    DFN1E1C0 \sr_10_[12]  (.D(\sr_9_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[12]_net_1 ));
    DFN1E1C0 \sr_26_[4]  (.D(\sr_25_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[4]_net_1 ));
    DFN1E1C0 \sr_47_[8]  (.D(\sr_46_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[8]_net_1 ));
    DFN1E1C0 \sr_44_[6]  (.D(\sr_43_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[6]_net_1 ));
    DFN1E1C0 \sr_42_[9]  (.D(\sr_41_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[9]_net_1 ));
    DFN1E1C0 \sr_63_[9]  (.D(\sr_62_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[9]));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \sr_10_[10]  (.D(\sr_9_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[10]_net_1 ));
    DFN1E1C0 \sr_2_[10]  (.D(sr_prev[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[10]_net_1 ));
    DFN1E1C0 \sr_13_[10]  (.D(\sr_12_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[10]_net_1 ));
    DFN1E1C0 \sr_57_[3]  (.D(\sr_56_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[3]_net_1 ));
    DFN1E1C0 \sr_27_[2]  (.D(\sr_26_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[2]_net_1 ));
    DFN1E1C0 \sr_40_[4]  (.D(\sr_39_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[4]_net_1 ));
    DFN1E1C0 \sr_30_[3]  (.D(\sr_29_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[3]_net_1 ));
    DFN1E1C0 \sr_50_[6]  (.D(\sr_49_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[6]_net_1 ));
    DFN1E1C0 \sr_27_[5]  (.D(\sr_26_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[5]_net_1 ));
    DFN1E1C0 \sr_46_[6]  (.D(\sr_45_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[6]_net_1 ));
    DFN1E1C0 \sr_38_[11]  (.D(\sr_37_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[11]_net_1 ));
    DFN1E1C0 \sr_17_[8]  (.D(\sr_16_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[8]_net_1 ));
    DFN1E1C0 \sr_20_[4]  (.D(\sr_19_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[4]_net_1 ));
    DFN1E1C0 \sr_0_[4]  (.D(cur_error[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[4]));
    DFN1E1C0 \sr_49_[11]  (.D(\sr_48_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[11]_net_1 ));
    DFN1E1C0 \sr_13_[9]  (.D(\sr_12_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[9]_net_1 ));
    DFN1E1C0 \sr_60_[6]  (.D(\sr_59_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[6]_net_1 ));
    DFN1E1C0 \sr_2_[7]  (.D(sr_prev[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[7]_net_1 ));
    DFN1E1C0 \sr_51_[1]  (.D(\sr_50_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[1]_net_1 ));
    DFN1E1C0 \sr_32_[0]  (.D(\sr_31_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[0]_net_1 ));
    DFN1E1C0 \sr_7_[2]  (.D(\sr_6_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[2]_net_1 ));
    DFN1E1C0 \sr_4_[11]  (.D(\sr_3_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[11]_net_1 ));
    DFN1E1C0 \sr_19_[2]  (.D(\sr_18_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[2]_net_1 ));
    DFN1E1C0 \sr_7_[8]  (.D(\sr_6_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[8]_net_1 ));
    DFN1E1C0 \sr_4_[5]  (.D(\sr_3_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[5]_net_1 ));
    DFN1E1C0 \sr_43_[0]  (.D(\sr_42_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[0]_net_1 ));
    DFN1E1C0 \sr_19_[0]  (.D(\sr_18_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[0]_net_1 ));
    DFN1E1C0 \sr_9_[10]  (.D(\sr_8_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[10]_net_1 ));
    DFN1E1C0 \sr_39_[8]  (.D(\sr_38_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[8]_net_1 ));
    DFN1E1C0 \sr_61_[1]  (.D(\sr_60_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[1]_net_1 ));
    DFN1E1C0 \sr_19_[10]  (.D(\sr_18_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[10]_net_1 ));
    DFN1E1C0 \sr_14_[1]  (.D(\sr_13_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[1]_net_1 ));
    DFN1E1C0 \sr_63_[3]  (.D(\sr_62_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[3]));
    DFN1E1C0 \sr_45_[7]  (.D(\sr_44_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[7]_net_1 ));
    DFN1E1C0 \sr_59_[5]  (.D(\sr_58_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[5]_net_1 ));
    DFN1E1C0 \sr_55_[7]  (.D(\sr_54_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[7]_net_1 ));
    DFN1E1C0 \sr_63_[12]  (.D(\sr_62_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[12]));
    DFN1E1C0 \sr_48_[1]  (.D(\sr_47_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[1]_net_1 ));
    DFN1E1C0 \sr_42_[12]  (.D(\sr_41_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[12]_net_1 ));
    DFN1E1C0 \sr_40_[6]  (.D(\sr_39_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[6]_net_1 ));
    DFN1E1C0 \sr_55_[8]  (.D(\sr_54_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[8]_net_1 ));
    DFN1E1C0 \sr_1_[4]  (.D(sr_new[4]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[4]));
    DFN1E1C0 \sr_34_[5]  (.D(\sr_33_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[5]_net_1 ));
    DFN1E1C0 \sr_6_[11]  (.D(\sr_5_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[11]_net_1 ));
    DFN1E1C0 \sr_11_[7]  (.D(\sr_10_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[7]_net_1 ));
    DFN1E1C0 \sr_34_[4]  (.D(\sr_33_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[4]_net_1 ));
    DFN1E1C0 \sr_16_[1]  (.D(\sr_15_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[1]_net_1 ));
    DFN1E1C0 \sr_29_[3]  (.D(\sr_28_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[3]_net_1 ));
    DFN1E1C0 \sr_17_[2]  (.D(\sr_16_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[2]_net_1 ));
    DFN1E1C0 \sr_39_[9]  (.D(\sr_38_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[9]_net_1 ));
    DFN1E1C0 \sr_3_[2]  (.D(\sr_2_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[2]_net_1 ));
    DFN1E1C0 \sr_46_[11]  (.D(\sr_45_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[11]_net_1 ));
    DFN1E1C0 \sr_3_[8]  (.D(\sr_2_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[8]_net_1 ));
    DFN1E1C0 \sr_33_[11]  (.D(\sr_32_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[11]_net_1 ));
    DFN1E1C0 \sr_17_[0]  (.D(\sr_16_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[0]_net_1 ));
    DFN1E1C0 \sr_37_[8]  (.D(\sr_36_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[8]_net_1 ));
    DFN1E1C0 \sr_15_[5]  (.D(\sr_14_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[5]_net_1 ));
    DFN1E1C0 \sr_11_[6]  (.D(\sr_10_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[6]_net_1 ));
    
endmodule


module controller_Z1_4_0(
       pwm_chg,
       sig_prev_0,
       sig_old_i_0_0,
       avg_done,
       N_46_1,
       pwm_rdy,
       sig_prev,
       sig_old_i_0,
       sum_rdy,
       deriv_enable,
       calc_avg,
       calc_int,
       pwm_enable,
       sum_enable,
       calc_error,
       avg_enable,
       int_enable,
       pwm_chg_0,
       avg_enable_0,
       n_rst_c,
       clk_c,
       avg_enable_1
    );
output pwm_chg;
input  sig_prev_0;
input  sig_old_i_0_0;
input  avg_done;
input  N_46_1;
input  pwm_rdy;
input  sig_prev;
input  sig_old_i_0;
input  sum_rdy;
output deriv_enable;
output calc_avg;
output calc_int;
output pwm_enable;
output sum_enable;
output calc_error;
output avg_enable;
output int_enable;
output pwm_chg_0;
output avg_enable_0;
input  n_rst_c;
input  clk_c;
output avg_enable_1;

    wire \state_RNII7JG[0]_net_1 , N_12, \state_1[5] , count_n14, 
        count_c13, \count[14]_net_1 , N_62, count_n13, count_c12, 
        \count[13]_net_1 , count_n12, count_c11, \count[12]_net_1 , 
        count_n15, count_31_0, N_95, count_c10, \count[11]_net_1 , 
        count_c9, \count[10]_net_1 , count_c8, \count[9]_net_1 , 
        count_c7, \count[8]_net_1 , count_c6, \count[7]_net_1 , 
        count_c5, \count[6]_net_1 , count_c4, \count[5]_net_1 , 
        count_c3, \count[4]_net_1 , count_c2, \count[3]_net_1 , 
        \count[1]_net_1 , \count[0]_net_1 , \count[2]_net_1 , 
        \state_ns_0_a2_9[0] , \state[10]_net_1 , N_33, 
        \state_ns_0_a2_8[0] , \state_ns_0_a2_6[0] , 
        \state_ns_0_a2_5[0] , \state_ns_0_a2_4[0] , N_272, 
        \state_ns_0_a2_1[0] , \state_ns_0_a2_0[0] , N_270, 
        \state[7]_net_1 , next_state_0_sqmuxa_1_1_a2_0_a2_0, 
        \state_ns_i_0_0[2] , un1_countlto15_13, un1_countlto15_5, 
        un1_countlto15_4, un1_countlto15_11, un1_countlto15_12, 
        un1_countlto15_1, un1_countlto15_0, un1_countlto15_9, 
        un1_countlto15_7, un1_countlto15_3, \count[15]_net_1 , 
        \state_RNO_0[5]_net_1 , N_24, N_274, N_273, \state[0]_net_1 , 
        N_23, N_26, next_state15_li, \state_RNIUI201[4]_net_1 , 
        count_n11, count_n10, count_n9, count_n2, count_n2_tz, 
        count_n3, count_n4, count_n5, count_n6, count_n7, count_n8, 
        \avg_count[0]_net_1 , \avg_count[1]_net_1 , \state_ns[1] , 
        \state_ns[0] , \state_ns[12] , \state[12]_net_1 , 
        \state_ns[7] , \state_ns[4] , \state[4]_net_1 , 
        \state_RNO_0[8] , \state_ns[10] , count_n1, N_267, counte, 
        \DWACT_ADD_CI_0_partial_sum[0] , I_10_0, 
        \DWACT_ADD_CI_0_TMP[0] , GND, VCC;
    
    DFN1E1C0 \count[5]  (.D(count_n5), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[5]_net_1 ));
    OA1A \state_RNO_0[0]  (.A(\state[10]_net_1 ), .B(N_33), .C(
        \state_ns_0_a2_8[0] ), .Y(\state_ns_0_a2_9[0] ));
    NOR2B \count_RNIK9SD1[7]  (.A(count_c6), .B(\count[7]_net_1 ), .Y(
        count_c7));
    DFN1E1C0 \count[1]  (.D(count_n1), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[1]_net_1 ));
    NOR2B \count_RNIQK481[6]  (.A(count_c5), .B(\count[6]_net_1 ), .Y(
        count_c6));
    NOR2 \count_RNILAFB[7]  (.A(\count[8]_net_1 ), .B(\count[7]_net_1 )
        , .Y(un1_countlto15_4));
    NOR2 \count_RNIFL9Q[13]  (.A(\count[14]_net_1 ), .B(
        \count[13]_net_1 ), .Y(un1_countlto15_1));
    DFN1E1C0 \count[10]  (.D(count_n10), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[10]_net_1 ));
    DFN1E1C0 \count[0]  (.D(N_267), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[0]_net_1 ));
    OR3C \state_RNO_9[0]  (.A(sig_old_i_0), .B(sig_prev), .C(
        \state[0]_net_1 ), .Y(N_270));
    DFN1C0 \state[13]  (.D(N_12), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_chg));
    NOR2B \count_RNIK5LJ2[11]  (.A(count_c10), .B(\count[11]_net_1 ), 
        .Y(count_c11));
    DFN1E1C0 \count[14]  (.D(count_n14), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[14]_net_1 ));
    OR2 \state_RNIDC64_0[4]  (.A(\state[12]_net_1 ), .B(
        \state[4]_net_1 ), .Y(N_272));
    DFN1C0 \state[7]  (.D(\state_ns[7] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[7]_net_1 ));
    NOR2B \count_RNI11D21[5]  (.A(count_c4), .B(\count[5]_net_1 ), .Y(
        count_c5));
    DFN1C0 \state[5]  (.D(\state_RNO_0[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_1[5] ));
    XA1B \count_RNO[7]  (.A(count_c6), .B(\count[7]_net_1 ), .C(N_62), 
        .Y(count_n7));
    AX1C \count_RNO[15]  (.A(count_c13), .B(count_31_0), .C(N_95), .Y(
        count_n15));
    NOR2 \count_RNI0ESI[9]  (.A(\count[10]_net_1 ), .B(
        \count[9]_net_1 ), .Y(un1_countlto15_3));
    AO1 \state_RNIALTT4[10]  (.A(sig_old_i_0_0), .B(sig_prev_0), .C(
        N_62), .Y(counte));
    DFN1C0 \state[4]  (.D(\state_ns[4] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[4]_net_1 ));
    NOR2A \count_RNO[2]  (.A(count_n2_tz), .B(N_62), .Y(count_n2));
    AO1A \state_RNO[7]  (.A(N_46_1), .B(\state[7]_net_1 ), .C(calc_int)
        , .Y(\state_ns[7] ));
    DFN1C0 \state_1[2]  (.D(\state_RNII7JG[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable_1));
    NOR3C \count_RNISB6H[2]  (.A(\count[1]_net_1 ), .B(
        \count[0]_net_1 ), .C(\count[2]_net_1 ), .Y(count_c2));
    NOR2A \state_RNO_0[5]  (.A(N_272), .B(\state[10]_net_1 ), .Y(N_24));
    DFN1C0 \state_0[2]  (.D(\state_RNII7JG[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable_0));
    XA1B \count_RNO[9]  (.A(count_c8), .B(\count[9]_net_1 ), .C(N_62), 
        .Y(count_n9));
    NOR2 \count_RNIH6FB[5]  (.A(\count[6]_net_1 ), .B(\count[5]_net_1 )
        , .Y(un1_countlto15_5));
    NOR2B \state_RNIUI201[4]  (.A(\state[4]_net_1 ), .B(avg_done), .Y(
        \state_RNIUI201[4]_net_1 ));
    DFN1C0 \state[6]  (.D(int_enable), .CLK(clk_c), .CLR(n_rst_c), .Q(
        calc_int));
    NOR3A \state_RNO_6[0]  (.A(N_270), .B(\state[7]_net_1 ), .C(
        sum_enable), .Y(\state_ns_0_a2_4[0] ));
    NOR2B \state_RNIPMAK[12]  (.A(\state[12]_net_1 ), .B(pwm_rdy), .Y(
        N_12));
    DFN1C0 \state[2]  (.D(\state_RNII7JG[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(avg_enable));
    VCC VCC_i (.Y(VCC));
    XOR2 un1_avg_count_1_I_10 (.A(\avg_count[1]_net_1 ), .B(
        \DWACT_ADD_CI_0_TMP[0] ), .Y(I_10_0));
    AOI1B \state_RNIA61H4[10]  (.A(un1_countlto15_13), .B(
        un1_countlto15_12), .C(next_state_0_sqmuxa_1_1_a2_0_a2_0), .Y(
        N_62));
    XA1B \count_RNO[4]  (.A(count_c3), .B(\count[4]_net_1 ), .C(N_62), 
        .Y(count_n4));
    DFN1C0 \state[3]  (.D(avg_enable), .CLK(clk_c), .CLR(n_rst_c), .Q(
        calc_avg));
    DFN1E1C0 \count[8]  (.D(count_n8), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[8]_net_1 ));
    XA1B \count_RNO[10]  (.A(count_c9), .B(\count[10]_net_1 ), .C(N_62)
        , .Y(count_n10));
    NOR2B \state_RNO[8]  (.A(\state[7]_net_1 ), .B(N_46_1), .Y(
        \state_RNO_0[8] ));
    NOR2 \count_RNIS9SI[15]  (.A(\count[15]_net_1 ), .B(
        \count[0]_net_1 ), .Y(un1_countlto15_0));
    NOR3B \state_RNO_1[0]  (.A(next_state15_li), .B(
        \state_RNIUI201[4]_net_1 ), .C(\state[10]_net_1 ), .Y(N_26));
    NOR3C \count_RNIMUBQ2[11]  (.A(un1_countlto15_1), .B(
        un1_countlto15_0), .C(un1_countlto15_9), .Y(un1_countlto15_12));
    NOR3A \count_RNIM0UM[3]  (.A(un1_countlto15_7), .B(
        \count[3]_net_1 ), .C(\count[4]_net_1 ), .Y(un1_countlto15_11));
    NOR2B \count_RNI9ELS[4]  (.A(count_c3), .B(\count[4]_net_1 ), .Y(
        count_c4));
    DFN1E1C0 \count[15]  (.D(count_n15), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[15]_net_1 ));
    XA1B \count_RNO[3]  (.A(count_c2), .B(\count[3]_net_1 ), .C(N_62), 
        .Y(count_n3));
    NOR2B \state_RNIOLO8[10]  (.A(\state[10]_net_1 ), .B(sum_rdy), .Y(
        next_state_0_sqmuxa_1_1_a2_0_a2_0));
    DFN1E1C0 \count[11]  (.D(count_n11), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[11]_net_1 ));
    DFN1C0 \state_0[13]  (.D(N_12), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_chg_0));
    XA1B \count_RNO[8]  (.A(count_c7), .B(\count[8]_net_1 ), .C(N_62), 
        .Y(count_n8));
    NOR3 \state_RNII7JG[0]  (.A(N_274), .B(\state_ns_i_0_0[2] ), .C(
        N_23), .Y(\state_RNII7JG[0]_net_1 ));
    AO1A \state_RNO[10]  (.A(sum_rdy), .B(\state[10]_net_1 ), .C(
        sum_enable), .Y(\state_ns[10] ));
    DFN1E1C0 \count[13]  (.D(count_n13), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[13]_net_1 ));
    XA1B \count_RNO[5]  (.A(count_c4), .B(\count[5]_net_1 ), .C(N_62), 
        .Y(count_n5));
    XA1B \count_RNO[1]  (.A(\count[1]_net_1 ), .B(\count[0]_net_1 ), 
        .C(N_62), .Y(count_n1));
    XA1B \count_RNO[11]  (.A(count_c10), .B(\count[11]_net_1 ), .C(
        N_62), .Y(count_n11));
    NOR2A \state_RNO_4[0]  (.A(\state_ns_0_a2_4[0] ), .B(N_272), .Y(
        \state_ns_0_a2_6[0] ));
    DFN1C0 \state[11]  (.D(N_62), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_enable));
    DFN1E1C0 \count[2]  (.D(count_n2), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[2]_net_1 ));
    NOR3A \count_RNIBV5D1[11]  (.A(un1_countlto15_3), .B(
        \count[11]_net_1 ), .C(\count[12]_net_1 ), .Y(un1_countlto15_9)
        );
    NOR2 \state_RNIOE85[0]  (.A(\state[0]_net_1 ), .B(N_272), .Y(N_23));
    NOR2B \count_RNIISTM[3]  (.A(count_c2), .B(\count[3]_net_1 ), .Y(
        count_c3));
    DFN1P0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .PRE(n_rst_c), 
        .Q(\state[0]_net_1 ));
    OR2B \state_RNIDC64[4]  (.A(\state[12]_net_1 ), .B(
        \state[4]_net_1 ), .Y(N_273));
    NOR3A \state_RNIKIC8[0]  (.A(N_273), .B(\state[10]_net_1 ), .C(
        \state[0]_net_1 ), .Y(N_274));
    DFN1C0 \state[12]  (.D(\state_ns[12] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[12]_net_1 ));
    NOR2A \count_RNO_1[15]  (.A(\count[15]_net_1 ), .B(N_62), .Y(N_95));
    GND GND_i (.Y(GND));
    DFN1E1C0 \count[9]  (.D(count_n9), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[9]_net_1 ));
    XA1B \count_RNO[6]  (.A(count_c5), .B(\count[6]_net_1 ), .C(N_62), 
        .Y(count_n6));
    XA1B \count_RNO[12]  (.A(count_c11), .B(\count[12]_net_1 ), .C(
        N_62), .Y(count_n12));
    NOR2 \count_RNO[0]  (.A(\count[0]_net_1 ), .B(N_62), .Y(N_267));
    NOR2B \count_RNIFVJJ1[8]  (.A(count_c7), .B(\count[8]_net_1 ), .Y(
        count_c8));
    AND2 un1_avg_count_1_I_1 (.A(\avg_count[0]_net_1 ), .B(
        \state_RNIUI201[4]_net_1 ), .Y(\DWACT_ADD_CI_0_TMP[0] ));
    XOR2 un1_avg_count_1_I_8 (.A(\avg_count[0]_net_1 ), .B(
        \state_RNIUI201[4]_net_1 ), .Y(\DWACT_ADD_CI_0_partial_sum[0] )
        );
    NOR2 \count_RNI9UEB[2]  (.A(\count[1]_net_1 ), .B(\count[2]_net_1 )
        , .Y(un1_countlto15_7));
    NOR2B \count_RNIBMBP1[9]  (.A(count_c8), .B(\count[9]_net_1 ), .Y(
        count_c9));
    NOR3B \state_RNO_5[0]  (.A(\state_ns_0_a2_1[0] ), .B(
        \state_ns_0_a2_0[0] ), .C(calc_error), .Y(\state_ns_0_a2_5[0] )
        );
    NOR3C \state_RNO_2[0]  (.A(un1_countlto15_12), .B(
        un1_countlto15_13), .C(sum_rdy), .Y(N_33));
    AO1A \state_RNO[4]  (.A(avg_done), .B(\state[4]_net_1 ), .C(
        calc_avg), .Y(\state_ns[4] ));
    NOR2B \count_RNI1PUD3[13]  (.A(count_c12), .B(\count[13]_net_1 ), 
        .Y(count_c13));
    DFN1E1C0 \count[6]  (.D(count_n6), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[6]_net_1 ));
    AO1A \state_RNO[12]  (.A(pwm_rdy), .B(\state[12]_net_1 ), .C(
        pwm_enable), .Y(\state_ns[12] ));
    DFN1C0 \state[10]  (.D(\state_ns[10] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[10]_net_1 ));
    NOR3C \count_RNISHSD1[3]  (.A(un1_countlto15_5), .B(
        un1_countlto15_4), .C(un1_countlto15_11), .Y(un1_countlto15_13)
        );
    DFN1E1C0 \count[3]  (.D(count_n3), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[3]_net_1 ));
    DFN1C0 \state[1]  (.D(\state_ns[1] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(calc_error));
    NOR2 \state_RNO_8[0]  (.A(calc_avg), .B(deriv_enable), .Y(
        \state_ns_0_a2_0[0] ));
    DFN1C0 \state[8]  (.D(\state_RNO_0[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(deriv_enable));
    OR3B \state_RNI66U2[7]  (.A(sig_old_i_0), .B(sig_prev), .C(
        \state[7]_net_1 ), .Y(\state_ns_i_0_0[2] ));
    AX1C \count_RNO_0[2]  (.A(\count[1]_net_1 ), .B(\count[0]_net_1 ), 
        .C(\count[2]_net_1 ), .Y(count_n2_tz));
    NOR3A \state_RNO[5]  (.A(calc_error), .B(\state[7]_net_1 ), .C(
        N_24), .Y(\state_RNO_0[5]_net_1 ));
    XA1B \count_RNO[14]  (.A(count_c13), .B(\count[14]_net_1 ), .C(
        N_62), .Y(count_n14));
    XA1B \count_RNO[13]  (.A(count_c12), .B(\count[13]_net_1 ), .C(
        N_62), .Y(count_n13));
    DFN1C0 \state[9]  (.D(deriv_enable), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(sum_enable));
    CLKINT \state_RNIG721[5]  (.A(\state_1[5] ), .Y(int_enable));
    NOR2B \count_RNIQUP03[12]  (.A(count_c11), .B(\count[12]_net_1 ), 
        .Y(count_c12));
    DFN1C0 \avg_count[0]  (.D(\DWACT_ADD_CI_0_partial_sum[0] ), .CLK(
        clk_c), .CLR(n_rst_c), .Q(\avg_count[0]_net_1 ));
    NOR2 \state_RNO_7[0]  (.A(pwm_enable), .B(calc_int), .Y(
        \state_ns_0_a2_1[0] ));
    AO1A \state_RNO[0]  (.A(int_enable), .B(\state_ns_0_a2_9[0] ), .C(
        N_26), .Y(\state_ns[0] ));
    DFN1C0 \avg_count[1]  (.D(I_10_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \avg_count[1]_net_1 ));
    OR2B \avg_count_RNI120A[1]  (.A(\avg_count[0]_net_1 ), .B(
        \avg_count[1]_net_1 ), .Y(next_state15_li));
    NOR2A \count_RNO_0[15]  (.A(\count[14]_net_1 ), .B(N_62), .Y(
        count_31_0));
    NOR3B \state_RNO_3[0]  (.A(\state_ns_0_a2_6[0] ), .B(
        \state_ns_0_a2_5[0] ), .C(avg_enable), .Y(\state_ns_0_a2_8[0] )
        );
    DFN1E1C0 \count[4]  (.D(count_n4), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[4]_net_1 ));
    NOR2B \count_RNIFDG62[10]  (.A(count_c9), .B(\count[10]_net_1 ), 
        .Y(count_c10));
    DFN1E1C0 \count[12]  (.D(count_n12), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[12]_net_1 ));
    NOR2A \state_RNO[1]  (.A(\state_RNIUI201[4]_net_1 ), .B(
        next_state15_li), .Y(\state_ns[1] ));
    DFN1E1C0 \count[7]  (.D(count_n7), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[7]_net_1 ));
    
endmodule


module sig_gen_2(
       primary_33_c,
       n_rst_c,
       clk_c,
       sig_old_i_0,
       sig_prev
    );
input  primary_33_c;
input  n_rst_c;
input  clk_c;
output sig_old_i_0;
output sig_prev;

    wire sig_prev_i, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(clk_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev_inst_1 (.D(primary_33_c), .CLK(clk_c), .CLR(
        n_rst_c), .Q(sig_prev));
    INV sig_old_RNO (.A(sig_prev), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module pid_sum_13s_4_0(
       integral_i,
       sr_new,
       integral,
       derivative_0,
       sr_new_0_0,
       sr_new_1_0,
       integral_0_0,
       integral_1_0,
       sum_39,
       sum_14,
       sum_19,
       sum_20,
       sum_22,
       sum_13,
       sum_18,
       sum_17,
       sum_21,
       sum_23,
       sum_16,
       sum_15,
       sum_12,
       sum_11,
       sum_6,
       sum_10,
       sum_9,
       sum_5,
       sum_8,
       sum_7,
       sum_4,
       sum_2_d0,
       sum_1_d0,
       sum_0_d0,
       sum_3,
       sum_0_0,
       sum_1_0,
       sum_2_0,
       sum_enable,
       sum_rdy,
       n_rst_c,
       clk_c
    );
input  [25:24] integral_i;
input  [12:0] sr_new;
input  [25:6] integral;
input  derivative_0;
input  sr_new_0_0;
input  sr_new_1_0;
input  integral_0_0;
input  integral_1_0;
output sum_39;
output sum_14;
output sum_19;
output sum_20;
output sum_22;
output sum_13;
output sum_18;
output sum_17;
output sum_21;
output sum_23;
output sum_16;
output sum_15;
output sum_12;
output sum_11;
output sum_6;
output sum_10;
output sum_9;
output sum_5;
output sum_8;
output sum_7;
output sum_4;
output sum_2_d0;
output sum_1_d0;
output sum_0_d0;
output sum_3;
output sum_0_0;
output sum_1_0;
output sum_2_0;
input  sum_enable;
output sum_rdy;
input  n_rst_c;
input  clk_c;

    wire \next_sum[39] , \state_RNIRSTG[6]_net_1 , \state_0[1]_net_1 , 
        \state_RNIGTM6[0]_net_1 , \state_2[2]_net_1 , 
        \state_1[2]_net_1 , \state_0[2]_net_1 , \state_0[3]_net_1 , 
        \state[6]_net_1 , N_416_0, \un1_next_sum_1_iv_0[26] , 
        \un1_next_sum_0_iv_0[25] , next_sum_1_sqmuxa, N_12, N_10, 
        \DWACT_FINC_E[0] , N_5, \DWACT_FINC_E[4] , N_2, 
        \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , N_25, N_23, 
        \DWACT_FINC_E_0[0] , N_18, \DWACT_FINC_E_0[4] , N_15, 
        \DWACT_FINC_E_0[7] , \DWACT_FINC_E_0[6] , N846, N778, N762, 
        N869, N785, I298_un1_Y, N882, N798, N814, I330_un1_Y, N838, 
        I338_un1_Y, N877, N1079, N881, I360_un1_Y, N666, N793, 
        I306_un1_Y, N770, N754, ADD_40x40_fast_I448_Y_0, 
        \sumreg[30]_net_1 , \un1_next_sum_1_iv[26] , 
        ADD_40x40_fast_I447_Y_0, \sumreg[29]_net_1 , 
        ADD_40x40_fast_I456_Y_0, \sumreg[38]_net_1 , 
        ADD_40x40_fast_I449_Y_0, \sumreg[31]_net_1 , 
        ADD_40x40_fast_I453_Y_0, \sumreg[35]_net_1 , 
        ADD_40x40_fast_I454_Y_0, \sumreg[36]_net_1 , 
        ADD_40x40_fast_I455_Y_0, \sumreg[37]_net_1 , 
        ADD_40x40_fast_I451_Y_0, \sumreg[33]_net_1 , 
        ADD_40x40_fast_I452_Y_0, \sumreg[34]_net_1 , 
        ADD_40x40_fast_I347_Y_0, N771, I284_un1_Y, 
        ADD_40x40_fast_I457_Y_0, ADD_40x40_fast_I446_Y_0, 
        \sumreg[28]_net_1 , ADD_40x40_fast_I450_Y_0, 
        \sumreg[32]_net_1 , ADD_40x40_fast_I379_Y_3, N756, 
        ADD_40x40_fast_I379_Y_2, N596, ADD_40x40_fast_I379_Y_0, N681, 
        ADD_40x40_fast_I382_Y_1, N777, ADD_40x40_fast_I382_Y_0, N679, 
        N687, ADD_40x40_fast_I381_Y_2, N760, N775, 
        ADD_40x40_fast_I381_Y_1, N600, N685, ADD_40x40_fast_I445_Y_0, 
        \sumreg[27]_net_1 , ADD_40x40_fast_I432_Y_0, 
        \un1_next_sum_iv_1[14] , \un1_next_sum_iv_2[14] , 
        ADD_40x40_fast_I380_Y_2, N758, N773, ADD_40x40_fast_I380_Y_1, 
        N598, N594, N683, ADD_40x40_fast_I347_un1_Y_0, N698, N690, 
        N788, ADD_40x40_fast_I437_Y_0, N_228_1, 
        \un1_next_sum_iv_0[19] , ADD_40x40_fast_I438_Y_0, 
        \un1_next_sum[20] , ADD_40x40_fast_I383_Y_1, N764, N779, 
        ADD_40x40_fast_I383_Y_0, N689, ADD_40x40_fast_I384_Y_1, N766, 
        N781, ADD_40x40_fast_I384_Y_0, N691, N684, 
        ADD_40x40_fast_I444_Y_0, \sumreg[26]_net_1 , 
        ADD_40x40_fast_I443_Y_0, \ireg_m[25] , 
        \un1_next_sum_0_iv_1[25] , \sumreg[25]_net_1 , 
        ADD_40x40_fast_I440_Y_0, \un1_next_sum[22] , 
        ADD_40x40_fast_I378_Y_3, N769, ADD_40x40_fast_I378_Y_2, 
        ADD_40x40_fast_I378_Y_0, N582, ADD_40x40_fast_I385_Y_2, 
        I280_un1_Y, ADD_40x40_fast_I385_Y_0, I385_un1_Y, N693, N686, 
        ADD_40x40_fast_I431_Y_0, \un1_next_sum[13] , 
        ADD_40x40_fast_I442_Y_0, \un1_next_sum_iv_0[24] , 
        \sumreg[24]_net_1 , ADD_40x40_fast_I436_Y_0, 
        \un1_next_sum_iv_1[18] , \un1_next_sum_iv_2[18] , 
        ADD_40x40_fast_I435_Y_0, \un1_next_sum[17] , 
        ADD_40x40_fast_I348_un1_Y_0, N790, N774, 
        ADD_40x40_fast_I439_Y_0, \un1_next_sum_iv_0[21] , 
        ADD_40x40_fast_I441_Y_0, \un1_next_sum_iv_0[23] , 
        ADD_40x40_fast_I434_Y_0, \un1_next_sum_iv_1[16] , 
        \un1_next_sum_iv_2[16] , ADD_40x40_fast_I433_Y_0, 
        \un1_next_sum_iv_1[15] , \un1_next_sum_iv_2[15] , 
        ADD_40x40_fast_I346_un1_Y_0, N786, ADD_40x40_fast_I430_Y_0, 
        \un1_next_sum[12] , ADD_40x40_fast_I349_un1_Y_0, N718, N710, 
        N776, ADD_40x40_fast_I429_Y_0, \un1_next_sum_iv_1[11] , 
        \un1_next_sum_iv_2[11] , ADD_40x40_fast_I380_un1_Y_0, N874, 
        N821, ADD_40x40_fast_I424_Y_0, \un1_next_sum[6] , 
        ADD_40x40_fast_I350_un1_Y_0, N794, ADD_40x40_fast_I428_Y_0, 
        \un1_next_sum_iv_1[10] , \un1_next_sum_iv_2[10] , 
        ADD_40x40_fast_I427_Y_0, \un1_next_sum_iv_1[9] , 
        \un1_next_sum_iv_2[9] , ADD_40x40_fast_I378_un1_Y_0, N802, 
        N817, ADD_40x40_fast_I382_un1_Y_0, N810, N743, 
        ADD_40x40_fast_I351_un1_Y_0, N796, N780, 
        ADD_40x40_fast_I423_Y_0, \un1_next_sum[5] , 
        ADD_40x40_fast_I426_Y_0, \un1_next_sum_iv_1[8] , 
        \un1_next_sum_iv_2[8] , ADD_40x40_fast_I384_un1_Y_0, 
        ADD_40x40_fast_I383_un1_Y_0, I116_un1_Y, N664, N880, 
        ADD_40x40_fast_I425_Y_0, \un1_next_sum[7] , 
        ADD_40x40_fast_I422_Y_0, \un1_next_sum_iv_0[4] , 
        ADD_40x40_fast_I420_Y_0, \un1_next_sum[0] , 
        ADD_40x40_fast_I419_Y_0, ADD_40x40_fast_I257_Y_1, N475, N472, 
        N661, ADD_40x40_fast_I201_Y_0, N601, N597, 
        ADD_40x40_fast_I197_Y_0, ADD_40x40_fast_I195_Y_0, 
        ADD_40x40_fast_I187_Y_0, ADD_22x22_fast_I179_Y_0, 
        \i_adj[21]_net_1 , \i_adj[19]_net_1 , ADD_22x22_fast_I126_Y_1, 
        N371, N378, ADD_22x22_fast_I126_Y_0, N335, N332, N331, 
        ADD_22x22_fast_I142_Y_0_1, ADD_22x22_fast_I142_Y_0_a3_0, N329, 
        ADD_22x22_fast_I142_Y_0_0, \i_adj[18]_net_1 , 
        \i_adj[20]_net_1 , N_14_1, ADD_22x22_fast_I172_Y_0, 
        \i_adj[14]_net_1 , \i_adj[12]_net_1 , 
        ADD_22x22_fast_I126_un1_Y_0, N379, ADD_22x22_fast_I175_Y_0, 
        \i_adj[17]_net_1 , \i_adj[15]_net_1 , 
        ADD_22x22_fast_I142_Y_0_a3_1, N330, ADD_40x40_fast_I418_Y_0, 
        ADD_22x22_fast_I177_Y_0, ADD_22x22_fast_I178_Y_0, 
        ADD_40x40_fast_I421_Y_0, ADD_22x22_fast_I130_Y_0, N386, 
        ADD_22x22_fast_I142_Y_0_o3_0_0, N337, N334, N333, 
        ADD_22x22_fast_I143_Y_3, ADD_22x22_fast_I143_un1_Y_0, N423, 
        ADD_22x22_fast_I143_Y_2, N367, N374, ADD_22x22_fast_I143_Y_1, 
        N328, ADD_22x22_fast_I143_Y_0, N314, ADD_22x22_fast_I144_Y_2, 
        ADD_22x22_fast_I144_un1_Y_0, N425, ADD_22x22_fast_I144_Y_1, 
        N369, N376, ADD_22x22_fast_I144_Y_0, \un1_next_sum_iv_0[20] , 
        \ireg[20]_net_1 , \state[3]_net_1 , \ireg[4]_net_1 , 
        \ireg[19]_net_1 , \ireg[21]_net_1 , \un1_next_sum_iv_0[5] , 
        \ireg[5]_net_1 , \ireg[23]_net_1 , \ireg[24]_net_1 , 
        \un1_next_sum_iv_0[22] , \ireg[22]_net_1 , 
        ADD_22x22_fast_I128_Y_0, N382, N375, ADD_22x22_fast_I170_Y_0, 
        \i_adj[10]_net_1 , ADD_22x22_fast_I169_Y_0, \i_adj[11]_net_1 , 
        \i_adj[9]_net_1 , \un1_next_sum_iv_2[6] , \un24_next_sum_m[6] , 
        next_sum_0_sqmuxa_1, \un3_next_sum_m[6] , 
        \un1_next_sum_iv_1[6] , \preg[6]_net_1 , next_sum_1_sqmuxa_2, 
        \ireg_m[6] , \un3_next_sum_m[16] , \un1_next_sum_iv_0[16] , 
        \ireg[16]_net_1 , \preg_m[16] , \preg[16]_net_1 , 
        next_sum_0_sqmuxa_2, \un3_next_sum_m[15] , 
        \un1_next_sum_iv_0[15] , \ireg[15]_net_1 , \preg_m[15] , 
        \preg[15]_net_1 , \un1_next_sum_iv_1[17] , \ireg[17]_net_1 , 
        \preg_m[17] , \un1_next_sum_iv_0[17] , \preg[17]_net_1 , 
        \ireg[14]_net_1 , next_sum_0_sqmuxa, \un1_next_sum_iv_0[14] , 
        \preg_m[14] , \preg[14]_net_1 , \un24_next_sum_m[8] , 
        \un3_next_sum_m[8] , \ireg[8]_net_1 , \preg_m[8] , 
        \un24_next_sum_m[10] , \un3_next_sum_m[10] , \preg[10]_net_1 , 
        \ireg_m[10] , \un24_next_sum_m[18] , \un3_next_sum_m[18] , 
        \ireg[18]_net_1 , \preg_m[18] , \un1_next_sum_iv_1[7] , 
        \preg[7]_net_1 , \ireg_m[7] , \un1_next_sum_iv_0[7] , 
        \un1_next_sum_iv_1[12] , \preg[12]_net_1 , \ireg_m[12] , 
        \un1_next_sum_iv_0[12] , \un24_next_sum_m[9] , 
        \un3_next_sum_m[9] , \ireg[9]_net_1 , \preg_m[9] , 
        \un24_next_sum_m[11] , \un3_next_sum_m[11] , \preg[11]_net_1 , 
        \ireg_m[11] , \un1_next_sum_iv_2[13] , \un24_next_sum_m[13] , 
        \un3_next_sum_m[13] , \un1_next_sum_iv_1[13] , 
        \preg[13]_net_1 , \ireg_m[13] , ADD_22x22_fast_I142_Y_0_a3_3_0, 
        N338, ADD_m8_i_1, ADD_m8_i_a4_0_1, N_232, \un3_next_sum_m[25] , 
        next_sum_1_sqmuxa_1, ADD_22x22_fast_I129_Y_0, N384, N377, 
        ADD_22x22_fast_I166_Y_0, \i_adj[8]_net_1 , \i_adj[6]_net_1 , 
        ADD_22x22_fast_I128_un1_Y_0, N383, ADD_22x22_fast_I131_Y_1, 
        ADD_22x22_fast_I131_Y_0, I131_un1_Y, N341, I72_un1_Y, 
        ADD_22x22_fast_I165_Y_0, \i_adj[7]_net_1 , \i_adj[5]_net_1 , 
        ADD_22x22_fast_I129_un1_Y_0, N385, N359, N266, 
        ADD_22x22_fast_I163_Y_0, \i_adj[3]_net_1 , N_9, 
        ADD_22x22_fast_I85_Y_0, \i_adj[4]_net_1 , \i_adj[2]_net_1 , 
        N270, ADD_m8_i_o4_1, ADD_m8_i_a4_1, N682, I352_un1_Y, N782, 
        N1103, N1055, I294_un1_Y, \un3_next_sum_m[12] , N1040, N1088, 
        I381_un1_Y, N876, N823, N844, N1027, I336_un1_Y, I383_un1_Y, 
        N848, N1035, N852, N883, N884, N1031, I340_un1_Y, N393, N354, 
        \next_ireg_3[15] , N424, I133_un1_Y, \next_ireg_3[7] , 
        \i_adj[1]_net_1 , N595, N599, I380_un1_Y, N1025, I334_un1_Y, 
        I349_un1_Y, N807, I317_un1_Y, N1046, I288_un1_Y, 
        \un3_next_sum_m[17] , \state[1]_net_1 , \next_ireg_3[25] , 
        N_12_0, \next_ireg_3[8] , \next_ireg_3[9] , N396, 
        \next_ireg_3[10] , N394, \next_ireg_3[16] , N422, I132_un1_Y, 
        \next_ireg_3[11] , N531, \next_ireg_3[13] , N525, 
        \next_ireg_3[19] , \i_adj[13]_net_1 , N507, \next_ireg_3[20] , 
        \i_adj[16]_net_1 , N504, \next_ireg_3[21] , N_17, 
        \next_ireg_3[22] , N498, \next_ireg_3[23] , I124_un1_Y, 
        \next_ireg_3[24] , I122_un1_Y, \next_ireg_3[18] , I130_un1_Y, 
        \next_ireg_3[17] , N513, \next_ireg_3[14] , N522, 
        \next_ireg_3[12] , N528, \un1_sumreg[11] , N809, I318_un1_Y, 
        \un1_sumreg[12] , \un1_sumreg[4] , \state[5]_net_1 , 
        \state[4]_net_1 , \un3_next_sum_m[7] , \un1_sumreg[2] , N1033, 
        I384_un1_Y, I342_un1_Y, N1029, I382_un1_Y, N1023, I332_un1_Y, 
        I379_un1_Y, N840, N872, N819, N1021, I378_un1_Y, N1058, 
        I296_un1_Y, N783, I353_un1_Y, N784, N800, N1106, N1052, 
        I292_un1_Y, I351_un1_Y, N1100, N1049, I290_un1_Y, I350_un1_Y, 
        N1043, I286_un1_Y, I348_un1_Y, N1091, N1037, I282_un1_Y, 
        I346_un1_Y, N1085, N680, N816, N734, \un1_sumreg[0] , 
        I106_un1_Y, N381, N389, N387, N740, N484, N481, 
        \inf_abs1_5[0] , \inf_abs1_5[1] , \inf_abs1_a_2[1] , 
        \inf_abs1_5[2] , \inf_abs1_a_2[2] , \inf_abs1_5[5] , 
        \inf_abs1_a_2[5] , N1070, N791, I304_un1_Y, I357_un1_Y, 
        \next_sum[20] , \inf_abs1_5[7] , \inf_abs1_a_2[7] , 
        \inf_abs1_5[10] , \inf_abs1_a_2[10] , \inf_abs2_5[1] , 
        \inf_abs2_a_0[1] , \inf_abs2_5[5] , \inf_abs2_a_0[5] , 
        \inf_abs2_5[12] , \inf_abs2_a_0[12] , \inf_abs2_5[13] , 
        \inf_abs2_a_0[13] , \inf_abs2_5[16] , \inf_abs2_a_0[16] , 
        \inf_abs2_5[17] , \inf_abs2_a_0[17] , \inf_abs2_5[18] , 
        \inf_abs2_a_0[18] , \inf_abs1_5[11] , \inf_abs1_a_2[11] , 
        \next_ireg_3[6] , \i_adj[0]_net_1 , \inf_abs2_5[0] , 
        \inf_abs2_5[2] , \inf_abs2_a_0[2] , \next_sum[0] , 
        \state[2]_net_1 , \next_sum[2] , \next_sum[4] , \next_sum[5] , 
        \next_sum[7] , \next_sum[8] , \next_sum[10] , \next_sum[11] , 
        \next_sum[12] , \next_sum[13] , \next_sum[16] , N1082, 
        \next_sum[18] , N1076, \next_sum[21] , N1067, \next_sum[22] , 
        N1064, \next_sum[23] , N1061, \next_sum[24] , \next_sum[27] , 
        \next_sum[29] , \next_sum[33] , \next_sum[35] , \next_sum[38] , 
        N276, N278, N282, N284, N288, N290, N291, N343, N347, N287, 
        N351, N281, N352, N355, N272, N275, N344, N348, N390, N391, 
        N356, N388, I114_un1_Y, N350, N346, N342, N297, N293, N296, 
        N345, N340, N300, N339, N299, N336, N315, N302, N303, N305, 
        N308, N309, N311, N312, N349, N353, N392, I115_un1_Y, N471, 
        N722, N641, N645, N725, N648, N644, N726, N649, I176_un1_Y, 
        N652, N729, N730, N653, N733, N656, N709, N702, N701, 
        I232_un1_Y, N717, N714, I240_un1_Y, N799, I252_un1_Y, 
        I184_un1_Y, N811, N812, N738, I256_un1_Y, N741, N815, 
        I259_un1_Y, I308_un1_Y, I312_un1_Y, I319_un1_Y, I359_un1_Y, 
        N795, I361_un1_Y, N657, N487, I236_un1_Y, N713, N636, N633, 
        N632, N519, N520, N721, N637, N514, N517, N706, N621, N538, 
        N541, N625, N629, N529, N526, N483, N486, N660, I164_un1_Y, 
        N513_0, N516, N640, N628, N525_0, N528_0, N624, N620, 
        I70_un1_Y, N540, N537, N495, N499, N498_0, N502, N505, N501, 
        N504_0, N496, N507_0, N510, N511, N642, N643, N647, N655, N490, 
        N658, N480, N723, N646, N724, N727, N650, N728, N651, N731, 
        N654, N732, N735, N736, I186_un1_Y, N662, N739, N704, N712, 
        I234_un1_Y, N719, N711, N720, I242_un1_Y, N801, N806, 
        I250_un1_Y, I254_un1_Y, N813, I314_un1_Y, N631, N630, N522_0, 
        N534, N535, N543, N544, N614, N546, N618, N619, N622, N623, 
        N634, N635, N612, N608, N611, N610, N692, N615, N695, N696, 
        N699, N700, N703, N626, N627, N705, N688, N707, N708, 
        I226_un1_Y, N787, I230_un1_Y, N715, N716, N797, N805, N808, 
        I300_un1_Y, I244_un1_Y, I302_un1_Y, N873, I310_un1_Y, 
        I315_un1_Y, I316_un1_Y, I320_un1_Y, I354_un1_Y, I355_un1_Y, 
        I358_un1_Y, \inf_abs2_5[3] , \inf_abs2_a_0[3] , 
        \inf_abs2_5[7] , \inf_abs2_a_0[7] , \inf_abs2_5[8] , 
        \inf_abs2_a_0[8] , \inf_abs2_5[19] , \inf_abs2_a_0[19] , 
        \inf_abs2_5[20] , \inf_abs2_a_0[20] , \inf_abs2_5[21] , 
        \inf_abs2_a_0[21] , \ireg[7]_net_1 , \preg[8]_net_1 , 
        \preg[9]_net_1 , \ireg[11]_net_1 , \ireg[13]_net_1 , 
        \preg[18]_net_1 , \state_ns[0] , \inf_abs2_5[14] , 
        \inf_abs2_a_0[14] , \inf_abs2_5[6] , \inf_abs2_a_0[6] , 
        \ireg[6]_net_1 , N489, N492, \next_sum[17] , \next_sum[6] , 
        N562, N559, N606, N565, N609, N603, N602, N694, \next_sum[28] , 
        \next_sum[37] , \next_sum[26] , \inf_abs1_5[12] , 
        \inf_abs1_a_2[12] , \inf_abs1_5[9] , \inf_abs1_a_2[9] , N357, 
        N269, I54_un1_Y, \next_sum[15] , \next_sum[34] , 
        \next_sum[32] , N604, \next_sum[1] , N1073, N532, N531_0, 
        \next_sum[36] , \next_sum[31] , \next_sum[19] , \next_sum[3] , 
        \inf_abs2_5[15] , \inf_abs2_a_0[15] , \inf_abs2_5[11] , 
        \inf_abs2_a_0[11] , \inf_abs2_5[10] , \inf_abs2_a_0[10] , 
        \inf_abs2_5[9] , \inf_abs2_a_0[9] , \inf_abs2_5[4] , 
        \inf_abs2_a_0[4] , \inf_abs1_5[6] , \inf_abs1_a_2[6] , 
        \next_sum[30] , \ireg[25]_net_1 , \ireg[12]_net_1 , 
        \ireg[10]_net_1 , \inf_abs1_5[8] , \inf_abs1_a_2[8] , 
        \inf_abs1_5[4] , \inf_abs1_a_2[4] , \inf_abs1_5[3] , 
        \inf_abs1_a_2[3] , N697, I212_un1_Y, N638, I144_un1_Y, N616, 
        N547, N613, I66_un1_Y, N550, I158_un1_Y, I166_un1_Y, 
        \next_sum[25] , \next_sum[14] , \next_sum[9] , 
        \p_adj[0]_net_1 , \p_adj[1]_net_1 , \p_adj[2]_net_1 , 
        \p_adj[3]_net_1 , \p_adj[4]_net_1 , \p_adj[5]_net_1 , 
        \p_adj[6]_net_1 , \p_adj[7]_net_1 , \p_adj[8]_net_1 , 
        \p_adj[9]_net_1 , \p_adj[10]_net_1 , \p_adj[11]_net_1 , 
        \p_adj[12]_net_1 , N_6, \DWACT_FINC_E[28] , \DWACT_FINC_E[13] , 
        \DWACT_FINC_E[15] , N_7, \DWACT_FINC_E[14] , N_8, 
        \DWACT_FINC_E[9] , \DWACT_FINC_E[12] , N_9_0, 
        \DWACT_FINC_E[10] , \DWACT_FINC_E[2] , \DWACT_FINC_E[5] , 
        N_10_0, \DWACT_FINC_E[11] , N_11, N_12_1, N_13, 
        \DWACT_FINC_E[8] , N_14, N_16, N_17_0, \DWACT_FINC_E[3] , N_19, 
        N_20, N_21, \DWACT_FINC_E[1] , N_22, N_24, N_3, 
        \DWACT_FINC_E_0[2] , \DWACT_FINC_E_0[5] , N_4, 
        \DWACT_FINC_E_0[3] , N_6_0, N_7_0, N_8_0, \DWACT_FINC_E_0[1] , 
        N_9_1, N_11_0, GND, VCC;
    
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I312_un1_Y (.A(N815), .B(N800), 
        .Y(I312_un1_Y));
    DFN1E1C0 \sumreg[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_39));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I77_Y (.A(N529), .B(N532), .Y(
        N627));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I19_G0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[19] ), .C(sum_19), .Y(N528_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I14_P0N (.A(
        \un1_next_sum_iv_1[14] ), .B(\un1_next_sum_iv_2[14] ), .C(
        sum_14), .Y(N514));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I46_Y (.A(\sumreg[34]_net_1 ), 
        .B(\sumreg[35]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N596)
        );
    XA1B \sumreg_RNO[10]  (.A(N1100), .B(ADD_40x40_fast_I428_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[10] ));
    MX2 \p_adj_RNO[2]  (.A(sr_new[2]), .B(\inf_abs1_a_2[2] ), .S(
        sr_new_1_0), .Y(\inf_abs1_5[2] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I336_un1_Y (.A(N791), .B(
        I304_un1_Y), .C(N844), .Y(I336_un1_Y));
    NOR2A \sumreg_RNO[11]  (.A(\un1_sumreg[11] ), .B(\state[2]_net_1 ), 
        .Y(\next_sum[11] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_0 (.A(N333), .B(N330), .C(
        N329), .Y(ADD_22x22_fast_I144_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I241_Y (.A(N726), .B(N718), .Y(
        N800));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I114_Y (.A(N471), .B(
        \un1_next_sum[0] ), .C(sum_1_d0), .Y(N664));
    DFN1E1C0 \i_adj[19]  (.D(\inf_abs2_5[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[19]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I113_Y (.A(N389), .B(N396), .C(
        N388), .Y(N525));
    DFN1E1C0 \sumreg[23]  (.D(\next_sum[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_23));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I290_un1_Y (.A(N793), .B(N778), 
        .Y(I290_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I128_un1_Y_0 (.A(N383), .B(N375)
        , .Y(ADD_22x22_fast_I128_un1_Y_0));
    NOR3B inf_abs1_a_2_I_19 (.A(\DWACT_FINC_E_0[2] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[6]), .Y(N_7_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I33_Y (.A(N303), .B(N300), .Y(
        N338));
    AND3 inf_abs2_a_0_I_30 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E_0[6] ));
    MX2 \i_adj_RNO[5]  (.A(integral[11]), .B(\inf_abs2_a_0[5] ), .S(
        integral_1_0), .Y(\inf_abs2_5[5] ));
    DFN1E1C0 \sumreg[38]  (.D(\next_sum[38] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(\sumreg[38]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I126_un1_Y_0 (.A(N371), .B(N379)
        , .Y(ADD_22x22_fast_I126_un1_Y_0));
    AO1A \ireg_RNI4DE12[14]  (.A(\ireg[14]_net_1 ), .B(
        next_sum_0_sqmuxa), .C(\un1_next_sum_iv_0[14] ), .Y(
        \un1_next_sum_iv_2[14] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I361_Y (.A(I361_un1_Y), .B(N883), 
        .Y(N1082));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I201_Y_0 (.A(N601), .B(N597), 
        .Y(ADD_40x40_fast_I201_Y_0));
    DFN1E1C0 \sumreg[5]  (.D(\next_sum[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_5));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I248_Y (.A(N733), .B(N726), .C(
        N725), .Y(N807));
    DFN1E1C0 \sumreg[20]  (.D(\next_sum[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_20));
    AO1 next_ireg_3_0_ADD_22x22_fast_I128_Y (.A(
        ADD_22x22_fast_I128_un1_Y_0), .B(N528), .C(
        ADD_22x22_fast_I128_Y_0), .Y(N504));
    NOR2 inf_abs2_a_0_I_57 (.A(integral[24]), .B(integral[25]), .Y(
        \DWACT_FINC_E[14] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I347_Y_0 (.A(N771), .B(
        I284_un1_Y), .Y(ADD_40x40_fast_I347_Y_0));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I52_Y (.A(\sumreg[32]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N602)
        );
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I199_Y (.A(N595), .B(N599), .C(
        N684), .Y(N758));
    DFN1E1C0 \sumreg[13]  (.D(\next_sum[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_13));
    NOR2A un1_sumreg_0_0_ADD_40x40_fast_I37_G0N (.A(\sumreg[37]_net_1 )
        , .B(\un1_next_sum_1_iv[26] ), .Y(N582));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I354_Y (.A(N785), .B(I298_un1_Y), 
        .C(I354_un1_Y), .Y(N1061));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I214_Y (.A(N699), .B(N692), .C(
        N691), .Y(N773));
    DFN1E1C0 \i_adj[2]  (.D(\inf_abs2_5[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[2]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I225_Y (.A(N702), .B(N710), .Y(
        N784));
    NOR3 \state_RNIALLC[6]  (.A(sum_rdy), .B(\state[6]_net_1 ), .C(
        \state_0[1]_net_1 ), .Y(N_416_0));
    NOR3A inf_abs1_a_2_I_13 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .C(
        sr_new[4]), .Y(N_9_1));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I436_Y_0 (.A(
        \un1_next_sum_iv_1[18] ), .B(\un1_next_sum_iv_2[18] ), .C(
        sum_18), .Y(ADD_40x40_fast_I436_Y_0));
    DFN1E1C0 \sumreg[27]  (.D(\next_sum[27] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[27]_net_1 ));
    DFN1E1C0 \sumreg[10]  (.D(\next_sum[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_10));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I381_Y_2 (.A(N760), .B(N775), .C(
        ADD_40x40_fast_I381_Y_1), .Y(ADD_40x40_fast_I381_Y_2));
    OR2 next_ireg_3_0_ADD_22x22_fast_I15_P0N (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(N312));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I444_Y_0 (.A(
        \sumreg[26]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I444_Y_0));
    XA1B \sumreg_RNO[22]  (.A(N1064), .B(ADD_40x40_fast_I440_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[22] ));
    NOR3B \preg_RNIFS18[9]  (.A(\state[5]_net_1 ), .B(\preg[9]_net_1 ), 
        .C(sr_new[12]), .Y(\preg_m[9] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I171_Y (.A(N643), .B(N647), .Y(
        N724));
    NOR2A \state_RNI170H_0[4]  (.A(\state[4]_net_1 ), .B(derivative_0), 
        .Y(next_sum_1_sqmuxa_1));
    OR2 next_ireg_3_0_ADD_22x22_fast_I11_P0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(N300));
    NOR2A \ireg_RNIAIG11_0[25]  (.A(next_sum_1_sqmuxa), .B(
        \ireg[25]_net_1 ), .Y(\un3_next_sum_m[25] ));
    AX1B un1_sumreg_0_0_ADD_40x40_fast_I443_Y_0 (.A(\ireg_m[25] ), .B(
        \un1_next_sum_0_iv_1[25] ), .C(\sumreg[25]_net_1 ), .Y(
        ADD_40x40_fast_I443_Y_0));
    XA1 \ireg_RNIML1B[5]  (.A(integral_0_0), .B(\ireg[5]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[5] ));
    AND2 inf_abs2_a_0_I_44 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E[9] ), .Y(\DWACT_FINC_E[10] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I18_P0N (.A(
        \un1_next_sum_iv_1[18] ), .B(\un1_next_sum_iv_2[18] ), .C(
        sum_18), .Y(N526));
    OR2 \ireg_RNI8FBP1[25]  (.A(\un1_next_sum_0_iv_0[25] ), .B(
        \un3_next_sum_m[25] ), .Y(\un1_next_sum_0_iv_1[25] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I306_un1_Y (.A(N809), .B(N794), 
        .Y(I306_un1_Y));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I166_Y (.A(I166_un1_Y), .B(N638), 
        .Y(N719));
    OA1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_0_0 (.A(
        \i_adj[18]_net_1 ), .B(\i_adj[20]_net_1 ), .C(N_9), .Y(
        ADD_22x22_fast_I142_Y_0_a3_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I10_P0N (.A(\i_adj[12]_net_1 ), 
        .B(\i_adj[10]_net_1 ), .Y(N297));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I168_Y (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[8]_net_1 ), .C(N522), .Y(\next_ireg_3[14] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I384_Y_1 (.A(N766), .B(N781), .C(
        ADD_40x40_fast_I384_Y_0), .Y(ADD_40x40_fast_I384_Y_1));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I10_G0N (.A(
        \un1_next_sum_iv_1[10] ), .B(\un1_next_sum_iv_2[10] ), .C(
        sum_10), .Y(N501));
    XNOR2 inf_abs1_a_2_I_28 (.A(sr_new[10]), .B(N_4), .Y(
        \inf_abs1_a_2[10] ));
    OR2 \state_RNIFSQA1[3]  (.A(N_228_1), .B(next_sum_0_sqmuxa), .Y(
        \un1_next_sum[0] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I18_G0N (.A(
        \un1_next_sum_iv_1[18] ), .B(\un1_next_sum_iv_2[18] ), .C(
        sum_18), .Y(N525_0));
    OR2 \preg_RNIPEM02[6]  (.A(\un1_next_sum_iv_2[6] ), .B(
        \un1_next_sum_iv_1[6] ), .Y(\un1_next_sum[6] ));
    AND2 un1_sumreg_0_0_ADD_40x40_fast_I338_un1_Y (.A(N877), .B(N846), 
        .Y(I338_un1_Y));
    DFN1E1C0 \p_adj[4]  (.D(\inf_abs1_5[4] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[4]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_2 (.A(
        ADD_22x22_fast_I144_un1_Y_0), .B(N425), .C(
        ADD_22x22_fast_I144_Y_1), .Y(ADD_22x22_fast_I144_Y_2));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I358_Y (.A(N793), .B(I306_un1_Y), 
        .C(I358_un1_Y), .Y(N1073));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I7_G0N (.A(\i_adj[9]_net_1 ), 
        .B(\i_adj[7]_net_1 ), .Y(N287));
    XNOR2 inf_abs2_a_0_I_20 (.A(integral[13]), .B(N_20), .Y(
        \inf_abs2_a_0[7] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I424_Y_0 (.A(sum_6), .B(
        \un1_next_sum[6] ), .Y(ADD_40x40_fast_I424_Y_0));
    DFN1E1C0 \sumreg[17]  (.D(\next_sum[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_17));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I257_Y_1 (.A(N475), .B(N472), 
        .C(N661), .Y(ADD_40x40_fast_I257_Y_1));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I321_Y (.A(N816), .B(
        \un1_next_sum[0] ), .C(N815), .Y(N1106));
    DFN1C0 \state[6]  (.D(\state[2]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[6]_net_1 ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I423_Y_0 (.A(sum_5), .B(
        \un1_next_sum[5] ), .Y(ADD_40x40_fast_I423_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y (.A(
        ADD_22x22_fast_I126_un1_Y_0), .B(N522), .C(
        ADD_22x22_fast_I126_Y_1), .Y(N498));
    AND3 inf_abs1_a_2_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[5] ), .Y(
        \DWACT_FINC_E[6] ));
    DFN1E1C0 \sumreg[35]  (.D(\next_sum[35] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(\sumreg[35]_net_1 ));
    MX2 \i_adj_RNO[13]  (.A(integral[19]), .B(\inf_abs2_a_0[13] ), .S(
        integral_0_0), .Y(\inf_abs2_5[13] ));
    DFN1E1C0 \sumreg[4]  (.D(\next_sum[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_4));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I166_Y_0 (.A(\i_adj[8]_net_1 ), 
        .B(\i_adj[6]_net_1 ), .Y(ADD_22x22_fast_I166_Y_0));
    XA1B \sumreg_RNO[38]  (.A(N1023), .B(ADD_40x40_fast_I456_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[38] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I160_Y (.A(N636), .B(N633), .C(
        N632), .Y(N713));
    NOR3B \ireg_RNI29KN[10]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[10]_net_1 ), .Y(\un3_next_sum_m[10] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I342_un1_Y (.A(N782), .B(N766), 
        .C(N881), .Y(I342_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I207_Y (.A(N684), .B(N692), .Y(
        N766));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I232_Y (.A(I232_un1_Y), .B(N709), 
        .Y(N791));
    NOR2 inf_abs2_a_0_I_6 (.A(integral[6]), .B(integral[7]), .Y(N_25));
    NOR3B inf_abs2_a_0_I_45 (.A(\DWACT_FINC_E[10] ), .B(
        \DWACT_FINC_E_0[6] ), .C(integral[21]), .Y(N_11));
    NOR3 inf_abs1_a_2_I_29 (.A(sr_new[7]), .B(sr_new[6]), .C(sr_new[8])
        , .Y(\DWACT_FINC_E_0[5] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I252_Y (.A(I252_un1_Y), .B(N729), 
        .Y(N811));
    MX2 \p_adj_RNO[1]  (.A(sr_new[1]), .B(\inf_abs1_a_2[1] ), .S(
        sr_new_1_0), .Y(\inf_abs1_5[1] ));
    AO1 \preg_RNIS1PA1[11]  (.A(\preg[11]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[11] ), .Y(
        \un1_next_sum_iv_1[11] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I382_un1_Y (.A(N778), .B(N762), 
        .C(ADD_40x40_fast_I382_un1_Y_0), .Y(I382_un1_Y));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I252_un1_Y (.A(N656), .B(
        I184_un1_Y), .C(N730), .Y(I252_un1_Y));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I30_Y (.A(N302), .B(
        \i_adj[15]_net_1 ), .C(\i_adj[13]_net_1 ), .Y(N335));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I124_un1_Y (.A(N377), .B(N369), 
        .C(N424), .Y(I124_un1_Y));
    AND2 un1_sumreg_0_0_ADD_40x40_fast_I330_un1_Y (.A(N869), .B(N838), 
        .Y(I330_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I237_Y (.A(N722), .B(N714), .Y(
        N796));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I176_un1_Y (.A(N652), .B(N649), 
        .Y(I176_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I12_G0N (.A(\i_adj[12]_net_1 ), 
        .B(\i_adj[14]_net_1 ), .Y(N302));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I422_Y (.A(
        ADD_40x40_fast_I422_Y_0), .B(N823), .Y(\un1_sumreg[4] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I11_G0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(N299));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I58_Y (.A(\sumreg[28]_net_1 ), 
        .B(\sumreg[29]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N608)
        );
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I257_Y (.A(
        ADD_40x40_fast_I257_Y_1), .B(N734), .Y(N816));
    AO1A \preg_RNIV0VV[17]  (.A(\preg[17]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[17] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I35_Y (.A(N297), .B(N300), .Y(
        N340));
    DFN1E1C0 \sumreg[7]  (.D(\next_sum[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_7));
    DFN1E1C0 \ireg[12]  (.D(\next_ireg_3[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[12]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I126_Y (.A(N602), .B(N598), .Y(
        N679));
    NOR2A inf_abs2_a_0_I_11 (.A(\DWACT_FINC_E_0[0] ), .B(integral[9]), 
        .Y(N_23));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I166_Y (.A(
        ADD_22x22_fast_I166_Y_0), .B(N528), .Y(\next_ireg_3[12] ));
    NOR3B \preg_RNIF0JE[18]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[18]_net_1 ), .Y(\un24_next_sum_m[18] ));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I38_Y (.A(N290), .B(
        \i_adj[11]_net_1 ), .C(\i_adj[9]_net_1 ), .Y(N343));
    XNOR2 inf_abs2_a_0_I_46 (.A(integral[22]), .B(N_11), .Y(
        \inf_abs2_a_0[16] ));
    XOR2 inf_abs1_a_2_I_5 (.A(sr_new[0]), .B(sr_new[1]), .Y(
        \inf_abs1_a_2[1] ));
    XNOR2 inf_abs1_a_2_I_23 (.A(sr_new[8]), .B(N_6_0), .Y(
        \inf_abs1_a_2[8] ));
    NOR3B \preg_RNISUL7[6]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[6]_net_1 ), .Y(\un24_next_sum_m[6] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I310_Y (.A(I310_un1_Y), .B(N797), 
        .Y(N881));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I308_un1_Y (.A(N811), .B(N796), 
        .Y(I308_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I169_Y (.A(N641), .B(N645), .Y(
        N722));
    DFN1C0 \state[2]  (.D(\state[1]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[2]_net_1 ));
    DFN1E1C0 \i_adj[15]  (.D(\inf_abs2_5[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[15]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I41_Y (.A(N291), .B(N288), .Y(
        N346));
    DFN1E1C0 \i_adj[20]  (.D(\inf_abs2_5[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[20]_net_1 ));
    XNOR2 inf_abs2_a_0_I_37 (.A(integral[19]), .B(N_14), .Y(
        \inf_abs2_a_0[13] ));
    MX2 \i_adj_RNO[12]  (.A(integral[18]), .B(\inf_abs2_a_0[12] ), .S(
        integral_0_0), .Y(\inf_abs2_5[12] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I53_Y (.A(\sumreg[32]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N603)
        );
    AO1 next_ireg_3_0_ADD_22x22_fast_I86_Y (.A(N356), .B(N359), .C(
        N355), .Y(N394));
    AX1D next_ireg_3_0_ADD_22x22_fast_I170_Y (.A(N422), .B(I132_un1_Y), 
        .C(ADD_22x22_fast_I170_Y_0), .Y(\next_ireg_3[16] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I379_un1_Y (.A(N840), .B(N872), 
        .C(N819), .Y(I379_un1_Y));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_1 (.A(N369), .B(N376), .C(
        ADD_22x22_fast_I144_Y_0), .Y(ADD_22x22_fast_I144_Y_1));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I4_P0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[4] ), .C(sum_4), .Y(N484));
    DFN1E1C0 \p_adj[10]  (.D(\inf_abs1_5[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[10]_net_1 ));
    AO1 \preg_RNIQVOA1[10]  (.A(\preg[10]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[10] ), .Y(
        \un1_next_sum_iv_1[10] ));
    DFN1E1C0 \p_adj[5]  (.D(\inf_abs1_5[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[5]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I164_Y (.A(I164_un1_Y), .B(N636), 
        .Y(N717));
    DFN1E1C0 \sumreg[36]  (.D(\next_sum[36] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(\sumreg[36]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I56_Y (.A(\sumreg[29]_net_1 ), 
        .B(\sumreg[30]_net_1 ), .C(\un1_next_sum_1_iv[26] ), .Y(N606));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I172_Y (.A(N648), .B(N645), .C(
        N644), .Y(N725));
    NOR2B \p_adj_RNO[12]  (.A(\inf_abs1_a_2[12] ), .B(sr_new[12]), .Y(
        \inf_abs1_5[12] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I300_un1_Y (.A(N721), .B(
        I244_un1_Y), .C(N788), .Y(I300_un1_Y));
    DFN1E1C0 \p_adj[0]  (.D(\inf_abs1_5[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[0]_net_1 ));
    AND3 inf_abs2_a_0_I_51 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[28] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I354_un1_Y (.A(N786), .B(N802), 
        .C(N817), .Y(I354_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I317_un1_Y (.A(N808), .B(N823), 
        .Y(I317_un1_Y));
    DFN1E1C0 \sumreg[9]  (.D(\next_sum[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_9));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I181_Y (.A(N657), .B(N653), .Y(
        N734));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I216_Y (.A(N701), .B(N694), .C(
        N693), .Y(N775));
    OA1 un1_sumreg_0_0_ADD_m8_i_a4 (.A(N_232), .B(ADD_m8_i_o4_1), .C(
        next_sum_0_sqmuxa), .Y(ADD_m8_i_a4_1));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I4_G0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[4] ), .C(sum_4), .Y(N483));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I129_Y (.A(N562), .B(N565), .C(
        N601), .Y(N682));
    NOR2B \preg_RNISNUE[15]  (.A(\preg[15]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[15] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I50_Y (.A(N272), .B(N276), .C(
        N275), .Y(N355));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I144_un1_Y_0 (.A(N377), .B(N369)
        , .C(N266), .Y(ADD_22x22_fast_I144_un1_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I34_Y (.A(N296), .B(N300), .C(
        N299), .Y(N339));
    DFN1E1C0 \sumreg[31]  (.D(\next_sum[31] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(\sumreg[31]_net_1 ));
    DFN1E1C0 \sumreg[2]  (.D(\next_sum[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_2_d0));
    DFN1E1C0 \i_adj[7]  (.D(\inf_abs2_5[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[7]_net_1 ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I383_Y (.A(
        ADD_40x40_fast_I383_Y_1), .B(I383_un1_Y), .C(I340_un1_Y), .Y(
        N1031));
    MX2 \i_adj_RNO[8]  (.A(integral[14]), .B(\inf_abs2_a_0[8] ), .S(
        integral_1_0), .Y(\inf_abs2_5[8] ));
    OR3 \preg_RNIDIK63[12]  (.A(\un1_next_sum_iv_0[12] ), .B(
        \un3_next_sum_m[12] ), .C(\un1_next_sum_iv_1[12] ), .Y(
        \un1_next_sum[12] ));
    AO1 \ireg_RNIBEEG1[18]  (.A(\ireg[18]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[18] ), .Y(
        \un1_next_sum_iv_1[18] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I9_P0N (.A(
        \un1_next_sum_iv_1[9] ), .B(\un1_next_sum_iv_2[9] ), .C(sum_9), 
        .Y(N499));
    NOR3A inf_abs2_a_0_I_27 (.A(\DWACT_FINC_E_0[4] ), .B(integral[15]), 
        .C(integral[14]), .Y(N_17_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I105_Y (.A(N487), .B(N490), .Y(
        N655));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I10_G0N (.A(\i_adj[12]_net_1 ), 
        .B(\i_adj[10]_net_1 ), .Y(N296));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I351_un1_Y_0 (.A(N796), .B(
        N780), .Y(ADD_40x40_fast_I351_un1_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I108_Y (.A(N390), .B(N383), .C(
        N382), .Y(N422));
    MX2 \p_adj_RNO[3]  (.A(sr_new[3]), .B(\inf_abs1_a_2[3] ), .S(
        sr_new_1_0), .Y(\inf_abs1_5[3] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I435_Y_0 (.A(sum_17), .B(
        \un1_next_sum[17] ), .Y(ADD_40x40_fast_I435_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I146_Y (.A(N622), .B(N619), .C(
        N618), .Y(N699));
    AND3 inf_abs2_a_0_I_48 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[11] ), .Y(N_10_0));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I197_Y_0 (.A(\sumreg[36]_net_1 )
        , .B(\sumreg[37]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(
        ADD_40x40_fast_I197_Y_0));
    DFN1E1C0 \preg[16]  (.D(\p_adj[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[16]_net_1 ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I135_Y (.A(N562), .B(N559), .C(
        N611), .Y(N688));
    DFN1E1C0 \preg[17]  (.D(\p_adj[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[17]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I9_G0N (.A(\i_adj[9]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(N293));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I155_Y (.A(N627), .B(N631), .Y(
        N708));
    OR3 \preg_RNICA7N1[11]  (.A(\un24_next_sum_m[11] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[11] ), .Y(
        \un1_next_sum_iv_2[11] ));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I122_un1_Y (.A(N375), .B(N367), 
        .C(N422), .Y(I122_un1_Y));
    OR2 next_ireg_3_0_ADD_22x22_fast_I12_P0N (.A(\i_adj[12]_net_1 ), 
        .B(\i_adj[14]_net_1 ), .Y(N303));
    OR2 next_ireg_3_0_ADD_22x22_fast_I5_P0N (.A(\i_adj[5]_net_1 ), .B(
        \i_adj[7]_net_1 ), .Y(N282));
    DFN1E1C0 \i_adj[8]  (.D(\inf_abs2_5[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[8]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I94_Y (.A(N501), .B(N505), .C(
        N504_0), .Y(N644));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I73_Y (.A(N346), .B(N342), .Y(
        N381));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I174_Y (.A(\i_adj[16]_net_1 ), 
        .B(\i_adj[14]_net_1 ), .C(N504), .Y(\next_ireg_3[20] ));
    DFN1E1C0 \i_adj[17]  (.D(\inf_abs2_5[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[17]_net_1 ));
    AO1A \preg_RNISTUV[14]  (.A(\preg[14]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[14] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I140_Y (.A(N616), .B(N613), .C(
        N612), .Y(N693));
    MX2 \i_adj_RNO[3]  (.A(integral[9]), .B(\inf_abs2_a_0[3] ), .S(
        integral_1_0), .Y(\inf_abs2_5[3] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I74_Y (.A(N531_0), .B(N535), .C(
        N534), .Y(N624));
    XNOR2 inf_abs2_a_0_I_49 (.A(integral[23]), .B(N_10_0), .Y(
        \inf_abs2_a_0[17] ));
    XNOR2 inf_abs2_a_0_I_12 (.A(integral[10]), .B(N_23), .Y(
        \inf_abs2_a_0[4] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I319_Y (.A(I319_un1_Y), .B(N811), 
        .Y(N1100));
    XA1B \sumreg_RNO[18]  (.A(N1076), .B(ADD_40x40_fast_I436_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[18] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I383_un1_Y_0 (.A(I116_un1_Y), .B(
        N664), .C(N880), .Y(ADD_40x40_fast_I383_un1_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I306_Y (.A(N793), .B(I306_un1_Y), 
        .Y(N877));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I224_Y (.A(N709), .B(N702), .C(
        N701), .Y(N783));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I383_Y_0 (.A(N681), .B(N689), .Y(
        ADD_40x40_fast_I383_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I17_G0N (.A(\un1_next_sum[17] )
        , .B(sum_17), .Y(N522_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I356_Y (.A(N874), .B(N821), .C(
        N873), .Y(N1067));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I239_Y (.A(N716), .B(N724), .Y(
        N798));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I259_Y (.A(N656), .B(I184_un1_Y), 
        .C(I259_un1_Y), .Y(N819));
    NOR2B \i_adj_RNO[21]  (.A(\inf_abs2_a_0[21] ), .B(integral[25]), 
        .Y(\inf_abs2_5[21] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I116_un1_Y (.A(N472), .B(
        \un1_next_sum[0] ), .Y(I116_un1_Y));
    DFN1E1C0 \sumreg[6]  (.D(\next_sum[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_6));
    DFN1E1C0 \sumreg[0]  (.D(\next_sum[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_0_d0));
    DFN1E1C0 \preg[15]  (.D(\p_adj[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[15]_net_1 ));
    DFN1E1C0 \i_adj[10]  (.D(\inf_abs2_5[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[10]_net_1 ));
    NOR3B \ireg_RNI8FKN[16]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[16]_net_1 ), .Y(\un3_next_sum_m[16] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I144_un1_Y (.A(N544), .B(N547), 
        .C(N620), .Y(I144_un1_Y));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I452_Y_0 (.A(
        \sumreg[34]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I452_Y_0));
    DFN1E1C0 \ireg[24]  (.D(\next_ireg_3[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[24]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I351_un1_Y (.A(
        ADD_40x40_fast_I351_un1_Y_0), .B(N1100), .Y(I351_un1_Y));
    XNOR2 inf_abs2_a_0_I_43 (.A(integral[21]), .B(N_12_1), .Y(
        \inf_abs2_a_0[15] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I69_Y (.A(N338), .B(N342), .Y(
        N377));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I385_Y (.A(N852), .B(N883), .C(
        ADD_40x40_fast_I385_Y_2), .Y(N1035));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I184_un1_Y (.A(N660), .B(N657), 
        .Y(I184_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I149_Y (.A(N621), .B(N625), .Y(
        N702));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I67_Y (.A(N336), .B(N340), .Y(
        N375));
    OR2 next_ireg_3_0_ADD_22x22_fast_I54_Y (.A(N269), .B(I54_un1_Y), 
        .Y(N359));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I378_Y_2 (.A(N594), .B(
        ADD_40x40_fast_I378_Y_0), .C(N679), .Y(ADD_40x40_fast_I378_Y_2)
        );
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I360_Y (.A(N881), .B(I360_un1_Y), 
        .Y(N1079));
    NOR2B \preg_RNIRMUE[14]  (.A(\preg[14]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[14] ));
    MX2 \p_adj_RNO[0]  (.A(sr_new[0]), .B(sr_new[0]), .S(sr_new_1_0), 
        .Y(\inf_abs1_5[0] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I384_Y_0 (.A(N691), .B(N684), .C(
        N683), .Y(ADD_40x40_fast_I384_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I182_Y (.A(N658), .B(N655), .C(
        N654), .Y(N735));
    AND3 inf_abs2_a_0_I_52 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[12] ), .Y(N_9_0));
    NOR3A inf_abs2_a_0_I_31 (.A(\DWACT_FINC_E_0[6] ), .B(integral[15]), 
        .C(integral[16]), .Y(N_16));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I232_un1_Y (.A(N717), .B(N710), 
        .Y(I232_un1_Y));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I163_Y (.A(N511), .B(N514), .C(
        N635), .Y(N716));
    AO1 next_ireg_3_0_ADD_22x22_fast_I110_Y (.A(N392), .B(N385), .C(
        N384), .Y(N424));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I197_Y (.A(N597), .B(
        ADD_40x40_fast_I197_Y_0), .C(N682), .Y(N756));
    DFN1E1C0 \i_adj[18]  (.D(\inf_abs2_5[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[18]_net_1 ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I91_Y (.A(sum_12), .B(
        \un1_next_sum[12] ), .C(N511), .Y(N641));
    AO1D un1_sumreg_0_0_ADD_40x40_fast_I25_P0N (.A(
        \un1_next_sum_0_iv_1[25] ), .B(\ireg_m[25] ), .C(
        \sumreg[25]_net_1 ), .Y(N547));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I144_Y (.A(I144_un1_Y), .B(N616), 
        .Y(N697));
    NOR3B \preg_RNIARIE[13]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[13]_net_1 ), .Y(\un24_next_sum_m[13] ));
    MX2 \i_adj_RNO[16]  (.A(integral[22]), .B(\inf_abs2_a_0[16] ), .S(
        integral_0_0), .Y(\inf_abs2_5[16] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I71_Y (.A(N538), .B(N541), .Y(
        N621));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I95_Y (.A(N502), .B(N505), .Y(
        N645));
    AO1 \ireg_RNIBOUS[9]  (.A(\ireg[9]_net_1 ), .B(next_sum_1_sqmuxa), 
        .C(\preg_m[9] ), .Y(\un1_next_sum_iv_1[9] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I319_un1_Y (.A(I116_un1_Y), .B(
        N664), .C(N812), .Y(I319_un1_Y));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I161_Y (.A(\i_adj[3]_net_1 ), .B(
        \i_adj[1]_net_1 ), .C(N266), .Y(\next_ireg_3[7] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I70_Y (.A(N343), .B(N340), .C(
        N339), .Y(N378));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I75_Y (.A(N532), .B(N535), .Y(
        N625));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I168_Y (.A(N644), .B(N641), .C(
        N640), .Y(N721));
    MX2 \p_adj_RNO[6]  (.A(sr_new[6]), .B(\inf_abs1_a_2[6] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[6] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I379_Y_3 (.A(N756), .B(N771), .C(
        ADD_40x40_fast_I379_Y_2), .Y(ADD_40x40_fast_I379_Y_3));
    OR3 \preg_RNIS4JD1[9]  (.A(\un24_next_sum_m[9] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[9] ), .Y(
        \un1_next_sum_iv_2[9] ));
    MX2 \i_adj_RNO[1]  (.A(integral[7]), .B(\inf_abs2_a_0[1] ), .S(
        integral_1_0), .Y(\inf_abs2_5[1] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I75_Y (.A(N344), .B(N348), .Y(
        N383));
    GND GND_i (.Y(GND));
    OR2 next_ireg_3_0_ADD_22x22_fast_I3_P0N (.A(\i_adj[5]_net_1 ), .B(
        \i_adj[3]_net_1 ), .Y(N276));
    OR2A un1_sumreg_0_0_ADD_40x40_fast_I31_P0N (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[31]_net_1 ), .Y(N565));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I143_Y_0 (.A(\i_adj[17]_net_1 ), 
        .B(\i_adj[19]_net_1 ), .C(N314), .Y(ADD_22x22_fast_I143_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I244_un1_Y (.A(N729), .B(N722), 
        .Y(I244_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I348_un1_Y_0 (.A(N790), .B(
        N774), .Y(ADD_40x40_fast_I348_un1_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I314_Y (.A(I314_un1_Y), .B(N801), 
        .Y(N1085));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I320_Y (.A(I320_un1_Y), .B(N813), 
        .Y(N1103));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I284_un1_Y (.A(N698), .B(N690), 
        .C(N787), .Y(I284_un1_Y));
    MX2 \p_adj_RNO[5]  (.A(sr_new[5]), .B(\inf_abs1_a_2[5] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[5] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I378_Y_3 (.A(N754), .B(N769), .C(
        ADD_40x40_fast_I378_Y_2), .Y(ADD_40x40_fast_I378_Y_3));
    DFN1C0 \state[5]  (.D(\state[4]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[5]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I78_Y (.A(N351), .B(N348), .C(
        N347), .Y(N386));
    NOR2 inf_abs2_a_0_I_21 (.A(integral[12]), .B(integral[13]), .Y(
        \DWACT_FINC_E[3] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I418_Y_0 (.A(sum_0_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I418_Y_0));
    NOR3B \preg_RNI7OIE[10]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[10]_net_1 ), .Y(\un24_next_sum_m[10] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I87_Y (.A(N514), .B(N517), .Y(
        N637));
    OA1 next_ireg_3_0_ADD_22x22_fast_I29_Y (.A(\i_adj[15]_net_1 ), .B(
        \i_adj[13]_net_1 ), .C(N309), .Y(N334));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I22_P0N (.A(\un1_next_sum[22] ), 
        .B(sum_22), .Y(N538));
    NOR3A inf_abs1_a_2_I_31 (.A(\DWACT_FINC_E[6] ), .B(sr_new[9]), .C(
        sr_new[10]), .Y(N_3));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I27_Y (.A(N309), .B(N312), .Y(
        N332));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I223_Y (.A(N700), .B(N708), .Y(
        N782));
    DFN1E1C0 \ireg[6]  (.D(\next_ireg_3[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[6]_net_1 ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I334_un1_Y (.A(N774), .B(N758), 
        .C(N873), .Y(I334_un1_Y));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I349_un1_Y_0 (.A(N718), .B(
        N710), .C(N776), .Y(ADD_40x40_fast_I349_un1_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I294_un1_Y (.A(N797), .B(N782), 
        .Y(I294_un1_Y));
    NOR3A \state_RNIJNKO[4]  (.A(integral[25]), .B(\state[5]_net_1 ), 
        .C(\state[4]_net_1 ), .Y(N_232));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I23_G0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[23] ), .C(sum_23), .Y(N540));
    DFN1E1C0 \preg[6]  (.D(\p_adj[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[6]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I36_Y (.A(N293), .B(N297), .C(
        N296), .Y(N341));
    OR2 \ireg_RNIKIS21[5]  (.A(\un1_next_sum_iv_0[5] ), .B(N_228_1), 
        .Y(\un1_next_sum[5] ));
    NOR2 inf_abs1_a_2_I_6 (.A(sr_new[0]), .B(sr_new[1]), .Y(N_12));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I1_G0N (.A(\i_adj[1]_net_1 ), 
        .B(\i_adj[3]_net_1 ), .Y(N269));
    OR2 next_ireg_3_0_ADD_22x22_fast_I114_Y (.A(I114_un1_Y), .B(N390), 
        .Y(N528));
    AO13 un1_sumreg_0_0_ADD_40x40_fast_I64_Y (.A(\sumreg[26]_net_1 ), 
        .B(N546), .C(\un1_next_sum_1_iv_0[26] ), .Y(N614));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I457_Y_0 (.A(sum_39), .B(
        \un1_next_sum_1_iv[26] ), .Y(ADD_40x40_fast_I457_Y_0));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I186_un1_Y (.A(N484), .B(N481), 
        .C(N662), .Y(I186_un1_Y));
    XA1B \sumreg_RNO[34]  (.A(N1031), .B(ADD_40x40_fast_I452_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[34] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I81_Y (.A(N354), .B(N350), .Y(
        N389));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I128_Y (.A(N600), .B(N604), .Y(
        N681));
    DFN1E1C0 \sumreg[29]  (.D(\next_sum[29] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[29]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I99_Y (.A(N496), .B(N499), .Y(
        N649));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I169_Y_0 (.A(\i_adj[11]_net_1 ), 
        .B(\i_adj[9]_net_1 ), .Y(ADD_22x22_fast_I169_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I226_Y (.A(I226_un1_Y), .B(N703), 
        .Y(N785));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I442_Y_0 (.A(N_228_1), .B(
        \un1_next_sum_iv_0[24] ), .C(\sumreg[24]_net_1 ), .Y(
        ADD_40x40_fast_I442_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I212_Y (.A(I212_un1_Y), .B(N689), 
        .Y(N771));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I79_Y (.A(N529), .B(N526), .Y(
        N629));
    NOR3B \ireg_RNI3AKN[11]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[11]_net_1 ), .Y(\un3_next_sum_m[11] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I167_Y (.A(N511), .B(N514), .C(
        N643), .Y(N720));
    NOR3 inf_abs1_a_2_I_10 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2])
        , .Y(\DWACT_FINC_E[0] ));
    DFN1C0 \state_0[3]  (.D(\state[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_0[3]_net_1 ));
    DFN1E1C0 \ireg[21]  (.D(\next_ireg_3[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[21]_net_1 ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I281_Y (.A(N694), .B(N686), .C(
        N784), .Y(N852));
    XNOR2 inf_abs2_a_0_I_32 (.A(integral[17]), .B(N_16), .Y(
        \inf_abs2_a_0[11] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I350_un1_Y_0 (.A(N794), .B(
        N778), .Y(ADD_40x40_fast_I350_un1_Y_0));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I430_Y_0 (.A(sum_12), .B(
        \un1_next_sum[12] ), .Y(ADD_40x40_fast_I430_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I217_Y (.A(N694), .B(N702), .Y(
        N776));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I378_un1_Y (.A(N770), .B(N754), 
        .C(ADD_40x40_fast_I378_un1_Y_0), .Y(I378_un1_Y));
    AND2 un1_sumreg_0_0_ADD_40x40_fast_I275_Y (.A(N778), .B(N762), .Y(
        N846));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I164_un1_Y (.A(N640), .B(N637), 
        .Y(I164_un1_Y));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I15_P0N (.A(
        \un1_next_sum_iv_1[15] ), .B(\un1_next_sum_iv_2[15] ), .C(
        sum_15), .Y(N517));
    XA1B \sumreg_RNO[27]  (.A(N1049), .B(ADD_40x40_fast_I445_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[27] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I74_Y (.A(N347), .B(N344), .C(
        N343), .Y(N382));
    DFN1E1C0 \sumreg[19]  (.D(\next_sum[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_19));
    NOR3B \ireg_RNIAHKN[18]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[18]_net_1 ), .Y(\un3_next_sum_m[18] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I422_Y_0 (.A(N_228_1), .B(
        \un1_next_sum_iv_0[4] ), .C(sum_4), .Y(ADD_40x40_fast_I422_Y_0)
        );
    DFN1E1C0 \sumreg[8]  (.D(\next_sum[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_8));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I353_un1_Y (.A(N784), .B(N800), 
        .C(N1106), .Y(I353_un1_Y));
    NOR3B \ireg_RNINN201[13]  (.A(\state[3]_net_1 ), .B(
        \ireg[13]_net_1 ), .C(integral_1_0), .Y(\ireg_m[13] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I349_un1_Y (.A(N807), .B(
        I317_un1_Y), .C(ADD_40x40_fast_I349_un1_Y_0), .Y(I349_un1_Y));
    DFN1E1C0 \sumreg[28]  (.D(\next_sum[28] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[28]_net_1 ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I179_Y_0 (.A(\i_adj[21]_net_1 ), 
        .B(\i_adj[19]_net_1 ), .Y(ADD_22x22_fast_I179_Y_0));
    AO1 \ireg_RNI7AEG1[16]  (.A(\ireg[16]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[16] ), .Y(
        \un1_next_sum_iv_1[16] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I304_un1_Y (.A(N718), .B(N710), 
        .C(N807), .Y(I304_un1_Y));
    NOR2A \sumreg_RNO[0]  (.A(\un1_sumreg[0] ), .B(\state[2]_net_1 ), 
        .Y(\next_sum[0] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I430_Y (.A(N807), .B(I317_un1_Y)
        , .C(ADD_40x40_fast_I430_Y_0), .Y(\un1_sumreg[12] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I256_un1_Y (.A(N741), .B(N734), 
        .Y(I256_un1_Y));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I451_Y_0 (.A(
        \sumreg[33]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I451_Y_0));
    AO1 un1_sumreg_0_0_ADD_m8_i_1 (.A(ADD_m8_i_a4_0_1), .B(N_232), .C(
        N_228_1), .Y(ADD_m8_i_1));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I143_Y (.A(N615), .B(N619), .Y(
        N696));
    NOR3B \preg_RNIV1M7[9]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[9]_net_1 ), .Y(\un24_next_sum_m[9] ));
    AO1 \preg_RNIHD1F1[13]  (.A(\preg[13]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[13] ), .Y(
        \un1_next_sum_iv_1[13] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_1_0 (.A(
        ADD_22x22_fast_I142_Y_0_a3_0), .B(N330), .Y(
        ADD_22x22_fast_I142_Y_0_a3_1));
    DFN1C0 \state_2[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_2[2]_net_1 ));
    DFN1E1C0 \sumreg[18]  (.D(\next_sum[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_18));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I380_Y_1 (.A(N598), .B(N594), .C(
        N683), .Y(ADD_40x40_fast_I380_Y_1));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I61_Y (.A(\sumreg[28]_net_1 ), 
        .B(\sumreg[27]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N611)
        );
    NOR2B next_ireg_3_0_ADD_22x22_fast_I6_G0N (.A(\i_adj[6]_net_1 ), 
        .B(\i_adj[8]_net_1 ), .Y(N284));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I162_Y (.A(\i_adj[4]_net_1 ), .B(
        \i_adj[2]_net_1 ), .C(N359), .Y(\next_ireg_3[8] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I21_P0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[21] ), .C(sum_21), .Y(N535));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I243_Y (.A(N720), .B(N728), .Y(
        N802));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I127_Y (.A(N603), .B(N599), .Y(
        N680));
    DFN1E1C0 \p_adj[3]  (.D(\inf_abs1_5[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[3]_net_1 ));
    DFN1E1C0 \ireg[10]  (.D(\next_ireg_3[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[10]_net_1 ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I49_Y (.A(\i_adj[6]_net_1 ), .B(
        \i_adj[4]_net_1 ), .C(N276), .Y(N354));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I65_Y (.A(N550), .B(N547), .Y(
        N615));
    OA1 next_ireg_3_0_ADD_22x22_fast_I47_Y (.A(\i_adj[6]_net_1 ), .B(
        \i_adj[4]_net_1 ), .C(N282), .Y(N352));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I101_Y (.A(sum_7), .B(
        \un1_next_sum[7] ), .C(N496), .Y(N651));
    AND3 inf_abs2_a_0_I_22 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_19));
    DFN1E1C0 \sumreg[1]  (.D(\next_sum[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_1_d0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I449_Y_0 (.A(
        \sumreg[31]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I449_Y_0));
    XA1B \sumreg_RNO[20]  (.A(N1070), .B(ADD_40x40_fast_I438_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[20] ));
    DFN1E1C0 \sumreg_0[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_0_0));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I47_Y (.A(\sumreg[35]_net_1 ), 
        .B(\sumreg[34]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N597)
        );
    XNOR2 inf_abs1_a_2_I_32 (.A(sr_new[11]), .B(N_3), .Y(
        \inf_abs1_a_2[11] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I187_Y_0 (.A(\un1_next_sum[0] ), 
        .B(sum_2_d0), .C(N475), .Y(ADD_40x40_fast_I187_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I148_Y (.A(N624), .B(N621), .C(
        N620), .Y(N701));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I165_Y (.A(
        ADD_22x22_fast_I165_Y_0), .B(N531), .Y(\next_ireg_3[11] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I13_G0N (.A(\un1_next_sum[13] )
        , .B(sum_13), .Y(N510));
    XA1B \sumreg_RNO[21]  (.A(N1067), .B(ADD_40x40_fast_I439_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[21] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_3_0 (.A(N334), .B(
        N338), .Y(ADD_22x22_fast_I142_Y_0_a3_3_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I250_un1_Y (.A(N735), .B(N728), 
        .Y(I250_un1_Y));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I131_Y (.A(N562), .B(N559), .C(
        N603), .Y(N684));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I303_Y (.A(N806), .B(N790), .Y(
        N874));
    XNOR2 inf_abs1_a_2_I_20 (.A(sr_new[7]), .B(N_7_0), .Y(
        \inf_abs1_a_2[7] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I438_Y_0 (.A(sum_20), .B(
        \un1_next_sum[20] ), .Y(ADD_40x40_fast_I438_Y_0));
    DFN1E1C0 \sumreg[25]  (.D(\next_sum[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[25]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I246_Y (.A(N731), .B(N724), .C(
        N723), .Y(N805));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I151_Y (.A(N627), .B(N623), .Y(
        N704));
    XA1 \ireg_RNILK1B[4]  (.A(integral_0_0), .B(\ireg[4]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[4] ));
    OR2 \preg_RNI1S863[13]  (.A(\un1_next_sum_iv_2[13] ), .B(
        \un1_next_sum_iv_1[13] ), .Y(\un1_next_sum[13] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I176_Y (.A(I176_un1_Y), .B(N648), 
        .Y(N729));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I347_Y (.A(
        ADD_40x40_fast_I347_un1_Y_0), .B(N1088), .C(
        ADD_40x40_fast_I347_Y_0), .Y(N1040));
    DFN1E1C0 \ireg[23]  (.D(\next_ireg_3[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[23]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I106_un1_Y (.A(N381), .B(N388), 
        .Y(I106_un1_Y));
    NOR2B \state_RNITLQ6[5]  (.A(\state[5]_net_1 ), .B(sr_new[12]), .Y(
        next_sum_0_sqmuxa_2));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I429_Y_0 (.A(
        \un1_next_sum_iv_1[11] ), .B(\un1_next_sum_iv_2[11] ), .C(
        sum_11), .Y(ADD_40x40_fast_I429_Y_0));
    OR2 un1_sumreg_0_0_ADD_m8_i (.A(ADD_m8_i_1), .B(ADD_m8_i_a4_1), .Y(
        N743));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I9_G0N (.A(
        \un1_next_sum_iv_1[9] ), .B(\un1_next_sum_iv_2[9] ), .C(sum_9), 
        .Y(N498_0));
    XA1B \state_RNI7GK5P9[2]  (.A(N1021), .B(ADD_40x40_fast_I457_Y_0), 
        .C(\state[2]_net_1 ), .Y(\next_sum[39] ));
    NOR3B \ireg_RNIPOSK[6]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[6]_net_1 ), .Y(\un3_next_sum_m[6] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I447_Y_0 (.A(
        \sumreg[29]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I447_Y_0));
    AO1 \ireg_RNI58EG1[15]  (.A(\ireg[15]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[15] ), .Y(
        \un1_next_sum_iv_1[15] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I353_Y (.A(I296_un1_Y), .B(N783), 
        .C(I353_un1_Y), .Y(N1058));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I316_un1_Y (.A(N806), .B(N821), 
        .Y(I316_un1_Y));
    AND3 inf_abs2_a_0_I_60 (.A(integral_i[24]), .B(integral_i[25]), .C(
        integral_i[25]), .Y(\DWACT_FINC_E[15] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I170_Y (.A(N646), .B(N643), .C(
        N642), .Y(N723));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I166_un1_Y (.A(N511), .B(N514), 
        .C(N642), .Y(I166_un1_Y));
    DFN1E1C0 \sumreg[15]  (.D(\next_sum[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_15));
    DFN1E1C0 \ireg[5]  (.D(\i_adj[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[5]_net_1 ));
    DFN1E1C0 \ireg[25]  (.D(\next_ireg_3[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[25]_net_1 ));
    AO1 \preg_RNIFB1F1[12]  (.A(\preg[12]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[12] ), .Y(
        \un1_next_sum_iv_1[12] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I16_P0N (.A(\i_adj[16]_net_1 ), 
        .B(\i_adj[18]_net_1 ), .Y(N315));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I5_G0N (.A(\un1_next_sum[5] ), 
        .B(sum_5), .Y(N486));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I427_Y_0 (.A(
        \un1_next_sum_iv_1[9] ), .B(\un1_next_sum_iv_2[9] ), .C(sum_9), 
        .Y(ADD_40x40_fast_I427_Y_0));
    NOR2B \ireg_RNIAIG11[25]  (.A(\ireg[25]_net_1 ), .B(
        next_sum_0_sqmuxa), .Y(\ireg_m[25] ));
    DFN1E1C0 \p_adj[9]  (.D(\inf_abs1_5[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[9]_net_1 ));
    XNOR2 inf_abs1_a_2_I_17 (.A(sr_new[6]), .B(N_8_0), .Y(
        \inf_abs1_a_2[6] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I163_Y (.A(
        ADD_22x22_fast_I163_Y_0), .B(N396), .Y(\next_ireg_3[9] ));
    MX2 \i_adj_RNO[14]  (.A(integral[20]), .B(\inf_abs2_a_0[14] ), .S(
        integral_0_0), .Y(\inf_abs2_5[14] ));
    OR2A un1_sumreg_0_0_ADD_40x40_fast_I30_P0N (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[30]_net_1 ), .Y(N562));
    NOR3B \ireg_RNIRQSK[8]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[8]_net_1 ), .Y(\un3_next_sum_m[8] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I69_Y (.A(N544), .B(N541), .Y(
        N619));
    XA1B \sumreg_RNO[14]  (.A(N1088), .B(ADD_40x40_fast_I432_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[14] ));
    XA1B \sumreg_RNO[35]  (.A(N1029), .B(ADD_40x40_fast_I453_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[35] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I349_Y (.A(I288_un1_Y), .B(N775), 
        .C(I349_un1_Y), .Y(N1046));
    DFN1C0 \state[4]  (.D(\state_0[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[4]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I147_Y (.A(N623), .B(N619), .Y(
        N700));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I8_G0N (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[8]_net_1 ), .Y(N290));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_0 (.A(\i_adj[18]_net_1 )
        , .B(\i_adj[20]_net_1 ), .C(N_14_1), .Y(
        ADD_22x22_fast_I142_Y_0_0));
    NOR2B \state_RNIHVVI[3]  (.A(\state[3]_net_1 ), .B(integral[25]), 
        .Y(next_sum_0_sqmuxa));
    DFN1E1C0 \sumreg[26]  (.D(\next_sum[26] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[26]_net_1 ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I441_Y_0 (.A(N_228_1), .B(
        \un1_next_sum_iv_0[23] ), .C(sum_23), .Y(
        ADD_40x40_fast_I441_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I179_Y (.A(N651), .B(N655), .Y(
        N732));
    XA1B \sumreg_RNO[7]  (.A(N817), .B(ADD_40x40_fast_I425_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[7] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I11_P0N (.A(
        \un1_next_sum_iv_1[11] ), .B(\un1_next_sum_iv_2[11] ), .C(
        sum_11), .Y(N505));
    AND2 un1_sumreg_0_0_ADD_40x40_fast_I267_Y (.A(N770), .B(N754), .Y(
        N838));
    AO1 next_ireg_3_0_ADD_22x22_fast_I128_Y_0 (.A(N382), .B(N375), .C(
        N374), .Y(ADD_22x22_fast_I128_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I90_Y (.A(N507_0), .B(N511), .C(
        N510), .Y(N640));
    DFN1E1C0 \ireg[17]  (.D(\next_ireg_3[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[17]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I316_Y (.A(I316_un1_Y), .B(N805), 
        .Y(N1091));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I305_Y (.A(N718), .B(N710), .C(
        N808), .Y(N876));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I381_Y (.A(
        ADD_40x40_fast_I381_Y_2), .B(I381_un1_Y), .C(I336_un1_Y), .Y(
        N1027));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I219_Y (.A(N704), .B(N696), .Y(
        N778));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I102_Y (.A(N489), .B(sum_7), .C(
        \un1_next_sum[7] ), .Y(N652));
    NOR3C un1_sumreg_0_0_ADD_m8_i_a4_0_1 (.A(sum_1_d0), .B(sum_0_d0), 
        .C(sum_2_d0), .Y(ADD_m8_i_a4_0_1));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I70_Y (.A(I70_un1_Y), .B(N540), 
        .Y(N620));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I21_G0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[21] ), .C(sum_21), .Y(N534));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I195_Y (.A(N595), .B(
        ADD_40x40_fast_I195_Y_0), .C(N680), .Y(N754));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I421_Y_0 (.A(sum_3), .B(N743), 
        .Y(ADD_40x40_fast_I421_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I318_un1_Y (.A(N810), .B(N743), 
        .Y(I318_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I174_Y (.A(N650), .B(N647), .C(
        N646), .Y(N727));
    DFN1E1C0 \sumreg[16]  (.D(\next_sum[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_16));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I16_G0N (.A(\i_adj[16]_net_1 ), 
        .B(\i_adj[18]_net_1 ), .Y(N314));
    XNOR2 inf_abs2_a_0_I_14 (.A(integral[11]), .B(N_22), .Y(
        \inf_abs2_a_0[5] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I355_Y (.A(N787), .B(I300_un1_Y), 
        .C(I355_un1_Y), .Y(N1064));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I132_Y (.A(N608), .B(N604), .Y(
        N685));
    NOR3B \ireg_RNI4BKN[12]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[12]_net_1 ), .Y(\un3_next_sum_m[12] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I2_G0N (.A(\i_adj[2]_net_1 ), 
        .B(\i_adj[4]_net_1 ), .Y(N272));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I152_Y (.A(N628), .B(N625), .C(
        N624), .Y(N705));
    MX2 \p_adj_RNO[8]  (.A(sr_new[8]), .B(\inf_abs1_a_2[8] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[8] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I3_P0N (.A(sum_3), .B(
        \un1_next_sum[0] ), .Y(N481));
    AO1 next_ireg_3_0_ADD_22x22_fast_I76_Y (.A(N349), .B(N346), .C(
        N345), .Y(N384));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I352_un1_Y (.A(N782), .B(N798), 
        .C(N1103), .Y(I352_un1_Y));
    DFN1E1C0 \sumreg[21]  (.D(\next_sum[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_21));
    MX2 \p_adj_RNO[7]  (.A(sr_new[7]), .B(\inf_abs1_a_2[7] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[7] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I84_Y (.A(N516), .B(N520), .C(
        N519), .Y(N634));
    AO1 next_ireg_3_0_ADD_22x22_fast_I42_Y (.A(N284), .B(N288), .C(
        N287), .Y(N347));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I222_Y (.A(N707), .B(N700), .C(
        N699), .Y(N781));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I315_un1_Y (.A(N730), .B(N722), 
        .C(N819), .Y(I315_un1_Y));
    XA1B \sumreg_RNO[36]  (.A(N1027), .B(ADD_40x40_fast_I454_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[36] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I1_P0N (.A(sum_1_d0), .B(
        \un1_next_sum[0] ), .Y(N475));
    NOR2B \preg_RNIUPUE[17]  (.A(\preg[17]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[17] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I158_un1_Y (.A(N634), .B(N631), 
        .Y(I158_un1_Y));
    OA1 next_ireg_3_0_ADD_22x22_fast_I31_Y (.A(\i_adj[15]_net_1 ), .B(
        \i_adj[13]_net_1 ), .C(N303), .Y(N336));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I70_un1_Y (.A(N537), .B(N541), 
        .Y(I70_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I380_un1_Y_0 (.A(N874), .B(
        N821), .Y(ADD_40x40_fast_I380_un1_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I310_un1_Y (.A(N813), .B(N798), 
        .Y(I310_un1_Y));
    AO1 next_ireg_3_0_ADD_22x22_fast_I129_Y (.A(
        ADD_22x22_fast_I129_un1_Y_0), .B(N531), .C(
        ADD_22x22_fast_I129_Y_0), .Y(N507));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I346_un1_Y (.A(
        ADD_40x40_fast_I346_un1_Y_0), .B(N1085), .Y(I346_un1_Y));
    DFN1E1C0 \p_adj[1]  (.D(\inf_abs1_5[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[1]_net_1 ));
    NOR3A inf_abs1_a_2_I_27 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .C(
        sr_new[9]), .Y(N_4));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I186_Y (.A(I186_un1_Y), .B(N658), 
        .Y(N739));
    NOR2 inf_abs2_a_0_I_15 (.A(integral[9]), .B(integral[10]), .Y(
        \DWACT_FINC_E[1] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I434_Y_0 (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(ADD_40x40_fast_I434_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I227_Y (.A(N704), .B(N712), .Y(
        N786));
    DFN1E1C0 \p_adj[7]  (.D(\inf_abs1_5[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[7]_net_1 ));
    DFN1E1C0 \sumreg[11]  (.D(\next_sum[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_11));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I433_Y_0 (.A(
        \un1_next_sum_iv_1[15] ), .B(\un1_next_sum_iv_2[15] ), .C(
        sum_15), .Y(ADD_40x40_fast_I433_Y_0));
    XA1B \sumreg_RNO[33]  (.A(N1033), .B(ADD_40x40_fast_I451_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[33] ));
    DFN1E1C0 \ireg[19]  (.D(\next_ireg_3[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[19]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I236_un1_Y (.A(N721), .B(N714), 
        .Y(I236_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I320_un1_Y (.A(N814), .B(N666), 
        .Y(I320_un1_Y));
    MX2 \i_adj_RNO[10]  (.A(integral[16]), .B(\inf_abs2_a_0[10] ), .S(
        integral_0_0), .Y(\inf_abs2_5[10] ));
    XNOR2 inf_abs2_a_0_I_40 (.A(integral[20]), .B(N_13), .Y(
        \inf_abs2_a_0[14] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I385_Y_0 (.A(N693), .B(N686), .C(
        N685), .Y(ADD_40x40_fast_I385_Y_0));
    AND3 inf_abs2_a_0_I_54 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E[9] ), .C(\DWACT_FINC_E[12] ), .Y(
        \DWACT_FINC_E[13] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I180_Y (.A(N656), .B(N653), .C(
        N652), .Y(N733));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I167_Y (.A(\i_adj[9]_net_1 ), .B(
        \i_adj[7]_net_1 ), .C(N525), .Y(\next_ireg_3[13] ));
    OR2 \ireg_RNIJJUN1[20]  (.A(\un1_next_sum_iv_0[20] ), .B(N_228_1), 
        .Y(\un1_next_sum[20] ));
    NOR3B \ireg_RNINM1B[6]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[6]_net_1 ), .C(integral_0_0), .Y(\ireg_m[6] ));
    DFN1C0 \state[1]  (.D(\state_RNIGTM6[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[1]_net_1 ));
    OR3 \preg_RNIQ2JD1[8]  (.A(\un24_next_sum_m[8] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[8] ), .Y(
        \un1_next_sum_iv_2[8] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I382_Y (.A(
        ADD_40x40_fast_I382_Y_1), .B(I382_un1_Y), .C(I338_un1_Y), .Y(
        N1029));
    MX2 \p_adj_RNO[10]  (.A(sr_new[10]), .B(\inf_abs1_a_2[10] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[10] ));
    DFN1E1C0 \ireg[22]  (.D(\next_ireg_3[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[22]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I20_P0N (.A(\un1_next_sum[20] ), 
        .B(sum_20), .Y(N532));
    AX1D next_ireg_3_0_ADD_22x22_fast_I169_Y (.A(N424), .B(I133_un1_Y), 
        .C(ADD_22x22_fast_I169_Y_0), .Y(\next_ireg_3[15] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I114_un1_Y (.A(N391), .B(N359), 
        .Y(I114_un1_Y));
    NOR3B inf_abs2_a_0_I_16 (.A(\DWACT_FINC_E[1] ), .B(
        \DWACT_FINC_E_0[0] ), .C(integral[11]), .Y(N_21));
    NOR2A \state_RNITLQ6_0[5]  (.A(\state[5]_net_1 ), .B(sr_new[12]), 
        .Y(next_sum_1_sqmuxa_2));
    NOR3B inf_abs2_a_0_I_55 (.A(\DWACT_FINC_E[13] ), .B(
        \DWACT_FINC_E[28] ), .C(integral[24]), .Y(N_8));
    DFN1E1C0 \preg[13]  (.D(\p_adj[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[13]_net_1 ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3 (.A(N_17), .B(
        ADD_22x22_fast_I142_Y_0_o3_0_0), .C(
        ADD_22x22_fast_I142_Y_0_a3_1), .Y(N_12_0));
    DFN1E1C0 \i_adj[6]  (.D(\inf_abs2_5[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[6]_net_1 ));
    DFN1E1C0 \i_adj[4]  (.D(\inf_abs2_5[4] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[4]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I63_Y (.A(N336), .B(N332), .Y(
        N371));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I81_Y (.A(sum_17), .B(
        \un1_next_sum[17] ), .C(N526), .Y(N631));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I379_Y_2 (.A(N596), .B(
        ADD_40x40_fast_I379_Y_0), .C(N681), .Y(ADD_40x40_fast_I379_Y_2)
        );
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I230_un1_Y (.A(N715), .B(N708), 
        .Y(I230_un1_Y));
    MX2 \i_adj_RNO[18]  (.A(integral[24]), .B(\inf_abs2_a_0[18] ), .S(
        integral_1_0), .Y(\inf_abs2_5[18] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I250_Y (.A(I250_un1_Y), .B(N727), 
        .Y(N809));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I456_Y_0 (.A(
        \sumreg[38]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I456_Y_0));
    NOR2A inf_abs1_a_2_I_11 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .Y(
        N_10));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I429_Y (.A(N809), .B(I318_un1_Y)
        , .C(ADD_40x40_fast_I429_Y_0), .Y(\un1_sumreg[11] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I348_Y (.A(I286_un1_Y), .B(N773), 
        .C(I348_un1_Y), .Y(N1043));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I165_Y (.A(N641), .B(N637), .Y(
        N718));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I381_Y_1 (.A(N596), .B(N600), .C(
        N685), .Y(ADD_40x40_fast_I381_Y_1));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I92_Y (.A(N504_0), .B(sum_12), 
        .C(\un1_next_sum[12] ), .Y(N642));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I348_un1_Y (.A(
        ADD_40x40_fast_I348_un1_Y_0), .B(N1091), .Y(I348_un1_Y));
    DFN1E1C0 \i_adj[9]  (.D(\inf_abs2_5[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[9]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I85_Y (.A(N520), .B(N517), .Y(
        N635));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I11_G0N (.A(
        \un1_next_sum_iv_1[11] ), .B(\un1_next_sum_iv_2[11] ), .C(
        sum_11), .Y(N504_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I201_Y (.A(
        ADD_40x40_fast_I201_Y_0), .B(N686), .Y(N760));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I72_Y (.A(N534), .B(N538), .C(
        N537), .Y(N622));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I0_S (.A(\i_adj[2]_net_1 ), .B(
        \i_adj[0]_net_1 ), .Y(\next_ireg_3[6] ));
    DFN1E1C0 \i_adj[3]  (.D(\inf_abs2_5[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[3]_net_1 ));
    XA1B \sumreg_RNO[15]  (.A(N1085), .B(ADD_40x40_fast_I433_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[15] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I242_Y (.A(I242_un1_Y), .B(N719), 
        .Y(N801));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y_1 (.A(N371), .B(N378), .C(
        ADD_22x22_fast_I126_Y_0), .Y(ADD_22x22_fast_I126_Y_1));
    OR2 next_ireg_3_0_ADD_22x22_fast_I14_P0N (.A(\i_adj[16]_net_1 ), 
        .B(\i_adj[14]_net_1 ), .Y(N309));
    OA1 next_ireg_3_0_ADD_22x22_fast_I51_Y (.A(\i_adj[4]_net_1 ), .B(
        \i_adj[2]_net_1 ), .C(N276), .Y(N356));
    AX1D next_ireg_3_0_ADD_22x22_fast_I178_Y (.A(I122_un1_Y), .B(
        ADD_22x22_fast_I143_Y_3), .C(ADD_22x22_fast_I178_Y_0), .Y(
        \next_ireg_3[24] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I231_Y (.A(N716), .B(N708), .Y(
        N790));
    XNOR2 inf_abs2_a_0_I_56 (.A(integral[25]), .B(N_8), .Y(
        \inf_abs2_a_0[19] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I87_Y (.A(I54_un1_Y), .B(N357), 
        .Y(N396));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I251_Y (.A(N736), .B(N728), .Y(
        N810));
    DFN1E1C0 \sumreg[34]  (.D(\next_sum[34] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(\sumreg[34]_net_1 ));
    XA1 \ireg_RNI9HG11[24]  (.A(integral[25]), .B(\ireg[24]_net_1 ), 
        .C(\state[3]_net_1 ), .Y(\un1_next_sum_iv_0[24] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I340_un1_Y (.A(N795), .B(
        I308_un1_Y), .C(N848), .Y(I340_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I247_Y (.A(N724), .B(N732), .Y(
        N806));
    DFN1C0 \state_0[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_0[2]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I60_Y (.A(\sumreg[28]_net_1 ), 
        .B(\sumreg[27]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N610)
        );
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I385_un1_Y (.A(N884), .B(
        \un1_next_sum[0] ), .C(N852), .Y(I385_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I173_Y (.A(N649), .B(N645), .Y(
        N726));
    DFN1E1C0 \ireg[7]  (.D(\next_ireg_3[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[7]_net_1 ));
    XA1B \sumreg_RNO[28]  (.A(N1046), .B(ADD_40x40_fast_I446_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[28] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I380_un1_Y (.A(N774), .B(N758), 
        .C(ADD_40x40_fast_I380_un1_Y_0), .Y(I380_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I238_Y (.A(N723), .B(N716), .C(
        N715), .Y(N797));
    XA1B \sumreg_RNO[3]  (.A(\un1_next_sum[0] ), .B(
        ADD_40x40_fast_I421_Y_0), .C(\state[2]_net_1 ), .Y(
        \next_sum[3] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I269_Y (.A(N698), .B(N690), .C(
        N756), .Y(N840));
    DFN1E1C0 \preg[7]  (.D(\p_adj[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[7]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I44_Y (.A(\sumreg[36]_net_1 ), 
        .B(\sumreg[35]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N594)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I258_Y (.A(N736), .B(N743), .C(
        N735), .Y(N817));
    OR2 next_ireg_3_0_ADD_22x22_fast_I131_Y (.A(
        ADD_22x22_fast_I131_Y_1), .B(I106_un1_Y), .Y(N513));
    DFN1E1C0 \ireg[16]  (.D(\next_ireg_3[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[16]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I273_Y (.A(N760), .B(N776), .Y(
        N844));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I195_Y_0 (.A(\sumreg[37]_net_1 )
        , .B(\sumreg[38]_net_1 ), .C(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I195_Y_0));
    XA1B \sumreg_RNO[32]  (.A(N1035), .B(ADD_40x40_fast_I450_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[32] ));
    DFN1E1C0 \preg[10]  (.D(\p_adj[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[10]_net_1 ));
    NOR3B \preg_RNIU0M7[8]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[8]_net_1 ), .Y(\un24_next_sum_m[8] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I163_Y_0 (.A(\i_adj[3]_net_1 ), 
        .B(\i_adj[5]_net_1 ), .Y(ADD_22x22_fast_I163_Y_0));
    DFN1E1C0 \preg[18]  (.D(\p_adj[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[18]_net_1 ));
    NOR3 \state_RNIRSTG[6]  (.A(sum_rdy), .B(\state[6]_net_1 ), .C(
        \state[1]_net_1 ), .Y(\state_RNIRSTG[6]_net_1 ));
    NOR3 inf_abs2_a_0_I_18 (.A(integral[10]), .B(integral[9]), .C(
        integral[11]), .Y(\DWACT_FINC_E[2] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I6_P0N (.A(\un1_next_sum[6] ), 
        .B(sum_6), .Y(N490));
    XA1B \sumreg_RNO[8]  (.A(N1106), .B(ADD_40x40_fast_I426_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[8] ));
    OR3 \preg_RNIGE7N1[13]  (.A(\un24_next_sum_m[13] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[13] ), .Y(
        \un1_next_sum_iv_2[13] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I131_Y_1 (.A(
        ADD_22x22_fast_I131_Y_0), .B(I131_un1_Y), .Y(
        ADD_22x22_fast_I131_Y_1));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I23_Y (.A(N315), .B(N_9), .Y(
        N328));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I384_un1_Y_0 (.A(N798), .B(
        N814), .C(N666), .Y(ADD_40x40_fast_I384_un1_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I178_Y (.A(N654), .B(N651), .C(
        N650), .Y(N731));
    NOR2B inf_abs2_a_0_I_34 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .Y(N_15));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I98_Y (.A(N495), .B(N499), .C(
        N498_0), .Y(N648));
    NOR2 inf_abs2_a_0_I_47 (.A(integral[21]), .B(integral[22]), .Y(
        \DWACT_FINC_E[11] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I10_P0N (.A(
        \un1_next_sum_iv_1[10] ), .B(\un1_next_sum_iv_2[10] ), .C(
        sum_10), .Y(N502));
    NOR2 inf_abs1_a_2_I_21 (.A(sr_new[6]), .B(sr_new[7]), .Y(
        \DWACT_FINC_E_0[3] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I5_G0N (.A(\i_adj[5]_net_1 ), 
        .B(\i_adj[7]_net_1 ), .Y(N281));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I176_Y (.A(\i_adj[16]_net_1 ), 
        .B(\i_adj[18]_net_1 ), .C(N498), .Y(\next_ireg_3[22] ));
    NOR3 inf_abs2_a_0_I_8 (.A(integral[7]), .B(integral[6]), .C(
        integral[8]), .Y(N_24));
    XA1B \sumreg_RNO[16]  (.A(N1082), .B(ADD_40x40_fast_I434_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[16] ));
    OR3 \preg_RNIA87N1[10]  (.A(\un24_next_sum_m[10] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[10] ), .Y(
        \un1_next_sum_iv_2[10] ));
    NOR3B inf_abs2_a_0_I_19 (.A(\DWACT_FINC_E[2] ), .B(
        \DWACT_FINC_E_0[0] ), .C(integral[12]), .Y(N_20));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I78_Y (.A(N525_0), .B(N529), .C(
        N528_0), .Y(N628));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I132_un1_Y (.A(N423), .B(N359), 
        .Y(I132_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I0_CO1 (.A(\i_adj[0]_net_1 ), 
        .B(\i_adj[2]_net_1 ), .Y(N266));
    OR2A un1_sumreg_0_0_ADD_40x40_fast_I26_P0N (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[26]_net_1 ), .Y(N550));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I229_Y (.A(N706), .B(N714), .Y(
        N788));
    XA1B \sumreg_RNO[13]  (.A(N1091), .B(ADD_40x40_fast_I431_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[13] ));
    OR3 \preg_RNIMUID1[6]  (.A(\un24_next_sum_m[6] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[6] ), .Y(
        \un1_next_sum_iv_2[6] ));
    XNOR2 inf_abs2_a_0_I_7 (.A(integral[8]), .B(N_25), .Y(
        \inf_abs2_a_0[2] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I133_un1_Y (.A(N425), .B(N266), 
        .Y(I133_un1_Y));
    XNOR2 inf_abs2_a_0_I_35 (.A(integral[18]), .B(N_15), .Y(
        \inf_abs2_a_0[12] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I1_P0N (.A(\i_adj[1]_net_1 ), .B(
        \i_adj[3]_net_1 ), .Y(N270));
    XOR2 inf_abs2_a_0_I_5 (.A(integral[6]), .B(integral[7]), .Y(
        \inf_abs2_a_0[1] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I357_un1_Y (.A(N876), .B(N823), 
        .Y(I357_un1_Y));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I332_un1_Y (.A(N787), .B(
        I300_un1_Y), .C(N840), .Y(I332_un1_Y));
    AND3 inf_abs2_a_0_I_61 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[15] ), .Y(N_6));
    XA1 \ireg_RNI8GG11[23]  (.A(integral[25]), .B(\ireg[23]_net_1 ), 
        .C(\state[3]_net_1 ), .Y(\un1_next_sum_iv_0[23] ));
    AND3 inf_abs2_a_0_I_58 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[14] ), .Y(N_7));
    OR3 \preg_RNIDD212[7]  (.A(\un1_next_sum_iv_0[7] ), .B(
        \un3_next_sum_m[7] ), .C(\un1_next_sum_iv_1[7] ), .Y(
        \un1_next_sum[7] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I111_Y (.A(sum_2_d0), .B(sum_3), 
        .C(\un1_next_sum[0] ), .Y(N661));
    XA1B \sumreg_RNO[19]  (.A(N1073), .B(ADD_40x40_fast_I437_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[19] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I68_Y (.A(N341), .B(N338), .C(
        N337), .Y(N376));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I16_G0N (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(N519));
    XNOR2 inf_abs1_a_2_I_12 (.A(sr_new[4]), .B(N_10), .Y(
        \inf_abs1_a_2[4] ));
    XA1 \ireg_RNILM301[20]  (.A(integral_1_0), .B(\ireg[20]_net_1 ), 
        .C(\state[3]_net_1 ), .Y(\un1_next_sum_iv_0[20] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I446_Y_0 (.A(
        \sumreg[28]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I446_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I109_Y (.A(N391), .B(N383), .Y(
        N423));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I93_Y (.A(sum_12), .B(
        \un1_next_sum[12] ), .C(N505), .Y(N643));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I212_un1_Y (.A(N697), .B(N690), 
        .Y(I212_un1_Y));
    DFN1E1C0 \p_adj[12]  (.D(\inf_abs1_5[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[12]_net_1 ));
    DFN1E1C0 \p_adj[2]  (.D(\inf_abs1_5[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[2]_net_1 ));
    MX2 \i_adj_RNO[9]  (.A(integral[15]), .B(\inf_abs2_a_0[9] ), .S(
        integral_1_0), .Y(\inf_abs2_5[9] ));
    DFN1E1C0 \ireg[18]  (.D(\next_ireg_3[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[18]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_1 (.A(N328), .B(N331), .C(
        ADD_22x22_fast_I143_Y_0), .Y(ADD_22x22_fast_I143_Y_1));
    NOR3A inf_abs2_a_0_I_13 (.A(\DWACT_FINC_E_0[0] ), .B(integral[9]), 
        .C(integral[10]), .Y(N_22));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I313_Y (.A(N816), .B(N800), .Y(
        N884));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I73_Y (.A(N535), .B(N538), .Y(
        N623));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_3 (.A(
        ADD_22x22_fast_I143_un1_Y_0), .B(N423), .C(
        ADD_22x22_fast_I143_Y_2), .Y(ADD_22x22_fast_I143_Y_3));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I45_Y (.A(\sumreg[36]_net_1 ), 
        .B(\sumreg[35]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N595)
        );
    DFN1E1C0 \ireg[9]  (.D(\next_ireg_3[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[9]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I382_Y_0 (.A(N679), .B(N687), .Y(
        ADD_40x40_fast_I382_Y_0));
    DFN1E1C0 \preg[14]  (.D(\p_adj[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[14]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I96_Y (.A(N498_0), .B(N502), .C(
        N501), .Y(N646));
    XNOR2 inf_abs2_a_0_I_59 (.A(integral[25]), .B(N_7), .Y(
        \inf_abs2_a_0[20] ));
    NOR2B \state_RNI170H[4]  (.A(derivative_0), .B(\state[4]_net_1 ), 
        .Y(next_sum_0_sqmuxa_1));
    XA1 \ireg_RNITT201[19]  (.A(integral_1_0), .B(\ireg[19]_net_1 ), 
        .C(\state[3]_net_1 ), .Y(\un1_next_sum_iv_0[19] ));
    AND3 inf_abs2_a_0_I_24 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E_0[4] ));
    DFN1E1C0 \preg[9]  (.D(\p_adj[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[9]_net_1 ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I426_Y_0 (.A(
        \un1_next_sum_iv_1[8] ), .B(\un1_next_sum_iv_2[8] ), .C(sum_8), 
        .Y(ADD_40x40_fast_I426_Y_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I379_Y (.A(I332_un1_Y), .B(
        ADD_40x40_fast_I379_Y_3), .C(I379_un1_Y), .Y(N1023));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I76_Y (.A(N528_0), .B(N532), .C(
        N531_0), .Y(N626));
    DFN1P0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .PRE(n_rst_c), 
        .Q(sum_rdy));
    AO1 \ireg_RNI9CEG1[17]  (.A(\ireg[17]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[17] ), .Y(
        \un1_next_sum_iv_1[17] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I205_Y (.A(N690), .B(N682), .Y(
        N764));
    NOR2B inf_abs1_a_2_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_2));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I177_Y (.A(N653), .B(N649), .Y(
        N730));
    NOR3B inf_abs2_a_0_I_36 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .C(integral[18]), .Y(N_14));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I8_G0N (.A(
        \un1_next_sum_iv_1[8] ), .B(\un1_next_sum_iv_2[8] ), .C(sum_8), 
        .Y(N495));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_3 (.A(
        ADD_22x22_fast_I142_Y_0_a3_3_0), .B(N513), .Y(N_17));
    XA1B \sumreg_RNO[6]  (.A(N819), .B(ADD_40x40_fast_I424_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[6] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I71_Y (.A(N340), .B(N344), .Y(
        N379));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I145_Y (.A(N544), .B(N547), .C(
        N621), .Y(N698));
    AO1A \state_RNO[0]  (.A(sum_enable), .B(sum_rdy), .C(
        \state[5]_net_1 ), .Y(\state_ns[0] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I62_Y (.A(\sumreg[27]_net_1 ), 
        .B(\sumreg[26]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N612)
        );
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I380_Y (.A(I380_un1_Y), .B(
        ADD_40x40_fast_I380_Y_2), .C(I334_un1_Y), .Y(N1025));
    NOR3B \ireg_RNI3DQR[10]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[10]_net_1 ), .C(integral_1_0), .Y(\ireg_m[10] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I235_Y (.A(N720), .B(N712), .Y(
        N794));
    NOR2A \state_RNIHVVI_0[3]  (.A(\state[3]_net_1 ), .B(integral[25]), 
        .Y(next_sum_1_sqmuxa));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I455_Y_0 (.A(
        \sumreg[37]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I455_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I255_Y (.A(N740), .B(N732), .Y(
        N814));
    AO1 next_ireg_3_0_ADD_22x22_fast_I82_Y (.A(N355), .B(N352), .C(
        N351), .Y(N390));
    NOR2A inf_abs2_a_0_I_25 (.A(\DWACT_FINC_E_0[4] ), .B(integral[14]), 
        .Y(N_18));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I183_Y (.A(N484), .B(N481), .C(
        N655), .Y(N736));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I254_un1_Y (.A(N739), .B(N732), 
        .Y(I254_un1_Y));
    DFN1E1C0 \ireg[8]  (.D(\next_ireg_3[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[8]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I302_un1_Y (.A(N805), .B(N790), 
        .Y(I302_un1_Y));
    AND2 un1_sumreg_0_0_ADD_40x40_fast_I360_un1_Y (.A(N666), .B(N882), 
        .Y(I360_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I25_Y (.A(N312), .B(N315), .Y(
        N330));
    OA1 next_ireg_3_0_ADD_22x22_fast_I43_Y (.A(\i_adj[8]_net_1 ), .B(
        \i_adj[6]_net_1 ), .C(N288), .Y(N348));
    XNOR2 inf_abs1_a_2_I_35 (.A(sr_new[12]), .B(N_2), .Y(
        \inf_abs1_a_2[12] ));
    DFN1E1C0 \preg[8]  (.D(\p_adj[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[8]_net_1 ));
    XNOR2 inf_abs2_a_0_I_53 (.A(integral[24]), .B(N_9_0), .Y(
        \inf_abs2_a_0[18] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I301_Y (.A(N730), .B(N722), .C(
        N788), .Y(N872));
    DFN1E1C0 \i_adj[14]  (.D(\inf_abs2_5[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[14]_net_1 ));
    OR2A un1_sumreg_0_0_ADD_40x40_fast_I29_P0N (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[29]_net_1 ), .Y(N559));
    DFN1E1C0 \sumreg[32]  (.D(\next_sum[32] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(\sumreg[32]_net_1 ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I346_Y (.A(I282_un1_Y), .B(N769), 
        .C(I346_un1_Y), .Y(N1037));
    AO1 next_ireg_3_0_ADD_22x22_fast_I28_Y (.A(N305), .B(N309), .C(
        N308), .Y(N333));
    NOR3A un1_sumreg_0_0_ADD_40x40_fast_I25_G0N (.A(\sumreg[25]_net_1 )
        , .B(\ireg_m[25] ), .C(\un1_next_sum_0_iv_1[25] ), .Y(N546));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I249_Y (.A(N726), .B(N734), .Y(
        N808));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I351_Y (.A(I292_un1_Y), .B(N779), 
        .C(I351_un1_Y), .Y(N1052));
    MX2 \i_adj_RNO[6]  (.A(integral[12]), .B(\inf_abs2_a_0[6] ), .S(
        integral_1_0), .Y(\inf_abs2_5[6] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I314_un1_Y (.A(N802), .B(N817), 
        .Y(I314_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I188_Y (.A(N664), .B(N661), .C(
        N660), .Y(N741));
    AND3 inf_abs1_a_2_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(N_6_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I16_P0N (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(N520));
    AO1A \preg_RNITUUV[15]  (.A(\preg[15]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[15] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I49_Y (.A(\sumreg[34]_net_1 ), 
        .B(\sumreg[33]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N599)
        );
    XNOR2 inf_abs2_a_0_I_26 (.A(integral[15]), .B(N_18), .Y(
        \inf_abs2_a_0[9] ));
    NOR2A \sumreg_RNO[12]  (.A(\un1_sumreg[12] ), .B(\state[2]_net_1 ), 
        .Y(\next_sum[12] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I54_Y (.A(\sumreg[31]_net_1 ), 
        .B(\sumreg[30]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N604)
        );
    NOR2B \preg_RNIVQUE[18]  (.A(\preg[18]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[18] ));
    NOR3B \ireg_RNI7EKN[15]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[15]_net_1 ), .Y(\un3_next_sum_m[15] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I315_Y (.A(N721), .B(I244_un1_Y), 
        .C(I315_un1_Y), .Y(N1088));
    XA1 \ireg_RNI7FG11[22]  (.A(integral[25]), .B(\ireg[22]_net_1 ), 
        .C(\state[3]_net_1 ), .Y(\un1_next_sum_iv_0[22] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I112_Y (.A(sum_1_d0), .B(
        sum_2_d0), .C(\un1_next_sum[0] ), .Y(N662));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I177_Y_0 (.A(\i_adj[19]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(ADD_22x22_fast_I177_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I106_Y (.A(N483), .B(N487), .C(
        N486), .Y(N656));
    OR2 \state_RNIFSQA1_1[3]  (.A(\un1_next_sum_0_iv_0[25] ), .B(
        next_sum_1_sqmuxa), .Y(\un1_next_sum_1_iv[26] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I7_G0N (.A(\un1_next_sum[7] ), 
        .B(sum_7), .Y(N492));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I242_un1_Y (.A(N727), .B(N720), 
        .Y(I242_un1_Y));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I164_Y (.A(\i_adj[4]_net_1 ), .B(
        \i_adj[6]_net_1 ), .C(N394), .Y(\next_ireg_3[10] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_1 (.A(
        ADD_22x22_fast_I142_Y_0_a3_0), .B(N329), .C(
        ADD_22x22_fast_I142_Y_0_0), .Y(ADD_22x22_fast_I142_Y_0_1));
    XNOR2 inf_abs2_a_0_I_62 (.A(integral[25]), .B(N_6), .Y(
        \inf_abs2_a_0[21] ));
    OR2 \state_RNIUSQN[5]  (.A(next_sum_0_sqmuxa_1), .B(
        next_sum_0_sqmuxa_2), .Y(N_228_1));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I419_Y_0 (.A(sum_1_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I419_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I68_Y (.A(N540), .B(N544), .C(
        N543), .Y(N618));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I22_G0N (.A(\un1_next_sum[22] )
        , .B(sum_22), .Y(N537));
    NOR2 inf_abs2_a_0_I_38 (.A(integral[18]), .B(integral[19]), .Y(
        \DWACT_FINC_E[8] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I380_Y_2 (.A(N758), .B(N773), .C(
        ADD_40x40_fast_I380_Y_1), .Y(ADD_40x40_fast_I380_Y_2));
    NOR3 inf_abs2_a_0_I_41 (.A(integral[19]), .B(integral[18]), .C(
        integral[20]), .Y(\DWACT_FINC_E[9] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I282_un1_Y (.A(N785), .B(N770), 
        .Y(I282_un1_Y));
    MX2 \p_adj_RNO[9]  (.A(sr_new[9]), .B(\inf_abs1_a_2[9] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[9] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I136_Y (.A(N612), .B(N608), .Y(
        N689));
    DFN1E1C0 \sumreg[33]  (.D(\next_sum[33] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(\sumreg[33]_net_1 ));
    NOR2A \sumreg_RNO[2]  (.A(\un1_sumreg[2] ), .B(\state[2]_net_1 ), 
        .Y(\next_sum[2] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I156_Y (.A(N632), .B(N629), .C(
        N628), .Y(N709));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I100_Y (.A(N492), .B(N496), .C(
        N495), .Y(N650));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I165_Y_0 (.A(\i_adj[7]_net_1 ), 
        .B(\i_adj[5]_net_1 ), .Y(ADD_22x22_fast_I165_Y_0));
    DFN1E1C0 \i_adj[12]  (.D(\inf_abs2_5[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[12]_net_1 ));
    NOR2B \i_adj_RNO[19]  (.A(\inf_abs2_a_0[19] ), .B(integral[25]), 
        .Y(\inf_abs2_5[19] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I359_un1_Y (.A(I116_un1_Y), .B(
        N664), .C(N880), .Y(I359_un1_Y));
    OA1 next_ireg_3_0_ADD_22x22_fast_I39_Y (.A(\i_adj[11]_net_1 ), .B(
        \i_adj[9]_net_1 ), .C(N291), .Y(N344));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I143_un1_Y_0 (.A(N375), .B(N367)
        , .C(N359), .Y(ADD_22x22_fast_I143_un1_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y_0 (.A(N335), .B(N332), .C(
        N331), .Y(ADD_22x22_fast_I126_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I14_G0N (.A(\i_adj[16]_net_1 ), 
        .B(\i_adj[14]_net_1 ), .Y(N308));
    DFN1E1C0 \sumreg[30]  (.D(\next_sum[30] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(\sumreg[30]_net_1 ));
    AND3 inf_abs2_a_0_I_39 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E_0[7] ), .C(\DWACT_FINC_E[8] ), .Y(N_13));
    AO1 next_ireg_3_0_ADD_22x22_fast_I24_Y (.A(N311), .B(N315), .C(
        N314), .Y(N329));
    OA1 next_ireg_3_0_ADD_22x22_fast_I37_Y (.A(\i_adj[11]_net_1 ), .B(
        \i_adj[9]_net_1 ), .C(N297), .Y(N342));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I302_Y (.A(N707), .B(I230_un1_Y), 
        .C(I302_un1_Y), .Y(N873));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I292_un1_Y (.A(N795), .B(N780), 
        .Y(I292_un1_Y));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I130_Y (.A(N606), .B(N602), .Y(
        N683));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I80_Y (.A(N522_0), .B(N526), .C(
        N525_0), .Y(N630));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I346_un1_Y_0 (.A(N786), .B(
        N770), .Y(ADD_40x40_fast_I346_un1_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I288_un1_Y (.A(N791), .B(N776), 
        .Y(I288_un1_Y));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I0_G0N (.A(N_228_1), .B(N_232), 
        .C(sum_0_d0), .Y(N471));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I150_Y (.A(N626), .B(N623), .C(
        N622), .Y(N703));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I161_Y (.A(N633), .B(N637), .Y(
        N714));
    AO1 next_ireg_3_0_ADD_22x22_fast_I40_Y (.A(N287), .B(N291), .C(
        N290), .Y(N345));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I172_Y_0 (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[12]_net_1 ), .Y(ADD_22x22_fast_I172_Y_0));
    OA1A un1_sumreg_0_0_ADD_40x40_fast_I63_Y (.A(
        \un1_next_sum_1_iv_0[26] ), .B(\sumreg[27]_net_1 ), .C(N550), 
        .Y(N613));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I420_Y (.A(I116_un1_Y), .B(N664)
        , .C(ADD_40x40_fast_I420_Y_0), .Y(\un1_sumreg[2] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I187_Y (.A(N484), .B(N481), .C(
        ADD_40x40_fast_I187_Y_0), .Y(N740));
    NOR2A \sumreg_RNO[4]  (.A(\un1_sumreg[4] ), .B(\state[2]_net_1 ), 
        .Y(\next_sum[4] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I352_Y (.A(I294_un1_Y), .B(N781), 
        .C(I352_un1_Y), .Y(N1055));
    XA1B \sumreg_RNO[5]  (.A(N821), .B(ADD_40x40_fast_I423_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[5] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I175_Y_0 (.A(\i_adj[17]_net_1 ), 
        .B(\i_adj[15]_net_1 ), .Y(ADD_22x22_fast_I175_Y_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I378_Y (.A(
        ADD_40x40_fast_I378_Y_3), .B(I378_un1_Y), .C(I330_un1_Y), .Y(
        N1021));
    OA1 next_ireg_3_0_ADD_22x22_fast_I45_Y (.A(\i_adj[8]_net_1 ), .B(
        \i_adj[6]_net_1 ), .C(N282), .Y(N350));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I171_Y (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .C(N513), .Y(\next_ireg_3[17] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_o3_0_0 (.A(N337), .B(
        N334), .C(N333), .Y(ADD_22x22_fast_I142_Y_0_o3_0_0));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I432_Y_0 (.A(
        \un1_next_sum_iv_1[14] ), .B(\un1_next_sum_iv_2[14] ), .C(
        sum_14), .Y(ADD_40x40_fast_I432_Y_0));
    DFN1E1C0 \sumreg[37]  (.D(\next_sum[37] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(\sumreg[37]_net_1 ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I51_Y (.A(\sumreg[33]_net_1 ), 
        .B(\sumreg[32]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N601)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I383_Y_1 (.A(N764), .B(N779), .C(
        ADD_40x40_fast_I383_Y_0), .Y(ADD_40x40_fast_I383_Y_1));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I23_P0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[23] ), .C(sum_23), .Y(N541));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_2 (.A(N367), .B(N374), .C(
        ADD_22x22_fast_I143_Y_1), .Y(ADD_22x22_fast_I143_Y_2));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I66_Y (.A(I66_un1_Y), .B(N546), 
        .Y(N616));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I445_Y_0 (.A(
        \sumreg[27]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I445_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I298_un1_Y (.A(N801), .B(N786), 
        .Y(I298_un1_Y));
    OR2 \preg_RNI4DJN1[15]  (.A(\un3_next_sum_m[15] ), .B(
        \un1_next_sum_iv_0[15] ), .Y(\un1_next_sum_iv_2[15] ));
    NOR3B \preg_RNI8PIE[11]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[11]_net_1 ), .Y(\un24_next_sum_m[11] ));
    XNOR2 inf_abs2_a_0_I_28 (.A(integral[16]), .B(N_17_0), .Y(
        \inf_abs2_a_0[10] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I19_P0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[19] ), .C(sum_19), .Y(N529));
    AO1 \preg_RNI3G3J[6]  (.A(\preg[6]_net_1 ), .B(next_sum_1_sqmuxa_2)
        , .C(\ireg_m[6] ), .Y(\un1_next_sum_iv_1[6] ));
    NOR3 inf_abs2_a_0_I_33 (.A(integral[16]), .B(integral[15]), .C(
        integral[17]), .Y(\DWACT_FINC_E_0[7] ));
    DFN1C0 \state_1[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_1[2]_net_1 ));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I48_Y (.A(N275), .B(
        \i_adj[6]_net_1 ), .C(\i_adj[4]_net_1 ), .Y(N353));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I3_G0N (.A(sum_3), .B(
        \un1_next_sum[0] ), .Y(N480));
    MX2 \i_adj_RNO[4]  (.A(integral[10]), .B(\inf_abs2_a_0[4] ), .S(
        integral_1_0), .Y(\inf_abs2_5[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I210_Y (.A(N695), .B(N688), .C(
        N687), .Y(N769));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I15_G0N (.A(
        \un1_next_sum_iv_1[15] ), .B(\un1_next_sum_iv_2[15] ), .C(
        sum_15), .Y(N516));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I425_Y_0 (.A(sum_7), .B(
        \un1_next_sum[7] ), .Y(ADD_40x40_fast_I425_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I139_Y (.A(N611), .B(N615), .Y(
        N692));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I384_un1_Y (.A(N782), .B(N766), 
        .C(ADD_40x40_fast_I384_un1_Y_0), .Y(I384_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I277_Y (.A(N764), .B(N780), .Y(
        N848));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I159_Y (.A(N635), .B(N631), .Y(
        N712));
    DFN1E1C0 \i_adj[13]  (.D(\inf_abs2_5[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[13]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I104_Y (.A(N486), .B(N490), .C(
        N489), .Y(N654));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I115_un1_Y (.A(N393), .B(N266), 
        .Y(I115_un1_Y));
    AO1A \preg_RNIUVUV[16]  (.A(\preg[16]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[16] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I54_un1_Y (.A(N270), .B(N266), 
        .Y(I54_un1_Y));
    NOR3 inf_abs2_a_0_I_29 (.A(integral[13]), .B(integral[12]), .C(
        integral[14]), .Y(\DWACT_FINC_E[5] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I130_Y_0 (.A(N386), .B(N379), .C(
        N378), .Y(ADD_22x22_fast_I130_Y_0));
    DFN1E1C0 \preg[12]  (.D(\p_adj[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[12]_net_1 ));
    MX2 \i_adj_RNO[2]  (.A(integral[8]), .B(\inf_abs2_a_0[2] ), .S(
        integral_1_0), .Y(\inf_abs2_5[2] ));
    DFN1E1C0 \i_adj[5]  (.D(\inf_abs2_5[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[5]_net_1 ));
    DFN1E1C0 \ireg[20]  (.D(\next_ireg_3[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[20]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I379_Y_0 (.A(\sumreg[37]_net_1 )
        , .B(\sumreg[36]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(
        ADD_40x40_fast_I379_Y_0));
    OR3 un1_sumreg_0_0_ADD_m8_i_o4_1 (.A(sum_2_d0), .B(sum_1_d0), .C(
        sum_0_d0), .Y(ADD_m8_i_o4_1));
    AO1A un1_sumreg_0_0_ADD_40x40_fast_I378_Y_0 (.A(
        \un1_next_sum_1_iv_0[26] ), .B(\sumreg[38]_net_1 ), .C(N582), 
        .Y(ADD_40x40_fast_I378_Y_0));
    AO1 \ireg_RNI9MUS[8]  (.A(\ireg[8]_net_1 ), .B(next_sum_1_sqmuxa), 
        .C(\preg_m[8] ), .Y(\un1_next_sum_iv_1[8] ));
    OR2 \state_RNIFSQA1_0[3]  (.A(\un1_next_sum_0_iv_0[25] ), .B(
        next_sum_1_sqmuxa), .Y(\un1_next_sum_1_iv_0[26] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I134_Y (.A(N610), .B(N606), .Y(
        N687));
    DFN1E1C0 \i_adj[0]  (.D(\inf_abs2_5[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[0]_net_1 ));
    DFN1E1C0 \p_adj[6]  (.D(\inf_abs1_5[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[6]_net_1 ));
    MX2 \p_adj_RNO[4]  (.A(sr_new[4]), .B(\inf_abs1_a_2[4] ), .S(
        sr_new_1_0), .Y(\inf_abs1_5[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I154_Y (.A(N630), .B(N627), .C(
        N626), .Y(N707));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I211_Y (.A(N688), .B(N696), .Y(
        N770));
    OR3 \preg_RNIHT183[17]  (.A(\un1_next_sum_iv_0[17] ), .B(
        \un3_next_sum_m[17] ), .C(\un1_next_sum_iv_1[17] ), .Y(
        \un1_next_sum[17] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I12_G0N (.A(\un1_next_sum[12] )
        , .B(sum_12), .Y(N507_0));
    XA1B \sumreg_RNO[24]  (.A(N1058), .B(ADD_40x40_fast_I442_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[24] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I59_Y (.A(N328), .B(N332), .Y(
        N367));
    MX2 \i_adj_RNO[0]  (.A(integral[6]), .B(integral[6]), .S(
        integral_1_0), .Y(\inf_abs2_5[0] ));
    AND3 inf_abs2_a_0_I_42 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E_0[7] ), .C(\DWACT_FINC_E[9] ), .Y(N_12_1));
    OR2 next_ireg_3_0_ADD_22x22_fast_I17_P0N_i_o3 (.A(
        \i_adj[19]_net_1 ), .B(\i_adj[17]_net_1 ), .Y(N_9));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I218_Y (.A(N703), .B(N696), .C(
        N695), .Y(N777));
    XNOR2 inf_abs2_a_0_I_23 (.A(integral[14]), .B(N_19), .Y(
        \inf_abs2_a_0[8] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I66_Y (.A(N339), .B(N336), .C(
        N335), .Y(N374));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I44_Y (.A(N281), .B(
        \i_adj[8]_net_1 ), .C(\i_adj[6]_net_1 ), .Y(N349));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I439_Y_0 (.A(N_228_1), .B(
        \un1_next_sum_iv_0[21] ), .C(sum_21), .Y(
        ADD_40x40_fast_I439_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I234_un1_Y (.A(N719), .B(N712), 
        .Y(I234_un1_Y));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I450_Y_0 (.A(
        \sumreg[32]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I450_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I234_Y (.A(I234_un1_Y), .B(N711), 
        .Y(N793));
    NOR3 inf_abs1_a_2_I_33 (.A(sr_new[10]), .B(sr_new[9]), .C(
        sr_new[11]), .Y(\DWACT_FINC_E[7] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I384_Y (.A(I384_un1_Y), .B(
        ADD_40x40_fast_I384_Y_1), .C(I342_un1_Y), .Y(N1033));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I254_Y (.A(I254_un1_Y), .B(N731), 
        .Y(N813));
    MX2 \i_adj_RNO[7]  (.A(integral[13]), .B(\inf_abs2_a_0[7] ), .S(
        integral_1_0), .Y(\inf_abs2_5[7] ));
    DFN1E1C0 \i_adj[21]  (.D(\inf_abs2_5[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[21]_net_1 ));
    XA1B \sumreg_RNO[9]  (.A(N1103), .B(ADD_40x40_fast_I427_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[9] ));
    OA1A un1_sumreg_0_0_ADD_40x40_fast_I59_Y (.A(
        \un1_next_sum_1_iv_0[26] ), .B(\sumreg[28]_net_1 ), .C(N559), 
        .Y(N609));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I162_Y (.A(N638), .B(N635), .C(
        N634), .Y(N715));
    DFN1E1C0 \ireg[14]  (.D(\next_ireg_3[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[14]_net_1 ));
    DFN1E1C0 \p_adj[11]  (.D(\inf_abs1_5[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[11]_net_1 ));
    XA1 \ireg_RNIMN301[21]  (.A(integral_1_0), .B(\ireg[21]_net_1 ), 
        .C(\state[3]_net_1 ), .Y(\un1_next_sum_iv_0[21] ));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I82_Y (.A(N519), .B(sum_17), .C(
        \un1_next_sum[17] ), .Y(N632));
    DFN1E1C0 \i_adj[16]  (.D(\inf_abs2_5[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[16]_net_1 ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I178_Y_0 (.A(\i_adj[20]_net_1 ), 
        .B(\i_adj[18]_net_1 ), .Y(ADD_22x22_fast_I178_Y_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I131_Y_0 (.A(N341), .B(I72_un1_Y), 
        .Y(ADD_22x22_fast_I131_Y_0));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I437_Y_0 (.A(N_228_1), .B(
        \un1_next_sum_iv_0[19] ), .C(sum_19), .Y(
        ADD_40x40_fast_I437_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I13_P0N (.A(\un1_next_sum[13] ), 
        .B(sum_13), .Y(N511));
    AO1 next_ireg_3_0_ADD_22x22_fast_I32_Y (.A(N299), .B(N303), .C(
        N302), .Y(N337));
    MX2 \i_adj_RNO[11]  (.A(integral[17]), .B(\inf_abs2_a_0[11] ), .S(
        integral_0_0), .Y(\inf_abs2_5[11] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I15_G0N (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(N311));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I385_Y_2 (.A(I280_un1_Y), .B(
        ADD_40x40_fast_I385_Y_0), .C(I385_un1_Y), .Y(
        ADD_40x40_fast_I385_Y_2));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I298_Y (.A(N785), .B(I298_un1_Y), 
        .Y(N869));
    DFN1E1C0 \ireg[4]  (.D(\i_adj[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[4]_net_1 ));
    MX2 \p_adj_RNO[11]  (.A(sr_new[11]), .B(\inf_abs1_a_2[11] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[11] ));
    AX1D next_ireg_3_0_ADD_22x22_fast_I172_Y (.A(I130_un1_Y), .B(
        ADD_22x22_fast_I130_Y_0), .C(ADD_22x22_fast_I172_Y_0), .Y(
        \next_ireg_3[18] ));
    XA1B \sumreg_RNO[37]  (.A(N1025), .B(ADD_40x40_fast_I455_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[37] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I381_un1_Y (.A(N876), .B(N823), 
        .C(N844), .Y(I381_un1_Y));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I141_Y (.A(N544), .B(N547), .C(
        N613), .Y(N694));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I83_Y (.A(N356), .B(N352), .Y(
        N391));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I72_un1_Y (.A(N345), .B(N342), 
        .Y(I72_un1_Y));
    AO1A \preg_RNIE12P[7]  (.A(\preg[7]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[7] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I111_Y (.A(N393), .B(N385), .Y(
        N425));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I175_Y (.A(N651), .B(N647), .Y(
        N728));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I378_un1_Y_0 (.A(N786), .B(
        N802), .C(N817), .Y(ADD_40x40_fast_I378_un1_Y_0));
    NOR2B \preg_RNITOUE[16]  (.A(\preg[16]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[16] ));
    DFN1E1C0 \sumreg[24]  (.D(\next_sum[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[24]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I26_Y (.A(N308), .B(N312), .C(
        N311), .Y(N331));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I24_G0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[24] ), .C(\sumreg[24]_net_1 ), .Y(N543));
    AX1D next_ireg_3_0_ADD_22x22_fast_I175_Y (.A(N_17), .B(
        ADD_22x22_fast_I142_Y_0_o3_0_0), .C(ADD_22x22_fast_I175_Y_0), 
        .Y(\next_ireg_3[21] ));
    NOR3B \ireg_RNI4EQR[11]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[11]_net_1 ), .C(integral_1_0), .Y(\ireg_m[11] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I431_Y_0 (.A(sum_13), .B(
        \un1_next_sum[13] ), .Y(ADD_40x40_fast_I431_Y_0));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I382_un1_Y_0 (.A(N794), .B(
        N810), .C(N743), .Y(ADD_40x40_fast_I382_un1_Y_0));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I103_Y (.A(sum_7), .B(
        \un1_next_sum[7] ), .C(N490), .Y(N653));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I259_un1_Y (.A(I116_un1_Y), .B(
        N664), .C(N738), .Y(I259_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I88_Y (.A(N510), .B(N514), .C(
        N513_0), .Y(N638));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I0_P0N (.A(N_228_1), .B(N_232), 
        .C(sum_0_d0), .Y(N472));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I260_Y (.A(N740), .B(N666), .C(
        N739), .Y(N821));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I8_P0N (.A(
        \un1_next_sum_iv_1[8] ), .B(\un1_next_sum_iv_2[8] ), .C(sum_8), 
        .Y(N496));
    MX2 \i_adj_RNO[15]  (.A(integral[21]), .B(\inf_abs2_a_0[15] ), .S(
        integral_0_0), .Y(\inf_abs2_5[15] ));
    OR2 \ireg_RNI5CBP1[22]  (.A(\un1_next_sum_iv_0[22] ), .B(N_228_1), 
        .Y(\un1_next_sum[22] ));
    DFN1E1C0 \sumreg[14]  (.D(\next_sum[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_14));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I350_Y (.A(I290_un1_Y), .B(N777), 
        .C(I350_un1_Y), .Y(N1049));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I203_Y (.A(N680), .B(N688), .Y(
        N762));
    NOR2B \i_adj_RNO[20]  (.A(\inf_abs2_a_0[20] ), .B(integral[25]), 
        .Y(\inf_abs2_5[20] ));
    XNOR2 inf_abs1_a_2_I_14 (.A(sr_new[5]), .B(N_9_1), .Y(
        \inf_abs1_a_2[5] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I170_Y_0 (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[12]_net_1 ), .Y(ADD_22x22_fast_I170_Y_0));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I133_Y (.A(N562), .B(N565), .C(
        N609), .Y(N686));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I215_Y (.A(N700), .B(N692), .Y(
        N774));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I153_Y (.A(N625), .B(N629), .Y(
        N706));
    NOR3B \ireg_RNI5CKN[13]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[13]_net_1 ), .Y(\un3_next_sum_m[13] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I79_Y (.A(N348), .B(N352), .Y(
        N387));
    XA1B \sumreg_RNO[30]  (.A(N1040), .B(ADD_40x40_fast_I448_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[30] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I77_Y (.A(N350), .B(N346), .Y(
        N385));
    XNOR2 inf_abs2_a_0_I_9 (.A(integral[9]), .B(N_24), .Y(
        \inf_abs2_a_0[3] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I226_un1_Y (.A(N711), .B(N704), 
        .Y(I226_un1_Y));
    XA1B \sumreg_RNO[31]  (.A(N1037), .B(ADD_40x40_fast_I449_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[31] ));
    NOR3 inf_abs2_a_0_I_10 (.A(integral[7]), .B(integral[6]), .C(
        integral[8]), .Y(\DWACT_FINC_E_0[0] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I440_Y_0 (.A(sum_22), .B(
        \un1_next_sum[22] ), .Y(ADD_40x40_fast_I440_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I253_Y (.A(N738), .B(N730), .Y(
        N812));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I52_Y (.A(N269), .B(
        \i_adj[4]_net_1 ), .C(\i_adj[2]_net_1 ), .Y(N357));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I108_Y (.A(N480), .B(N484), .C(
        N483), .Y(N658));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I261_Y (.A(N741), .B(I116_un1_Y), 
        .Y(N823));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I173_Y (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[15]_net_1 ), .C(N507), .Y(\next_ireg_3[19] ));
    OR2 \preg_RNI6FJN1[16]  (.A(\un3_next_sum_m[16] ), .B(
        \un1_next_sum_iv_0[16] ), .Y(\un1_next_sum_iv_2[16] ));
    NOR3B \ireg_RNIMM201[12]  (.A(\state[3]_net_1 ), .B(
        \ireg[12]_net_1 ), .C(integral_1_0), .Y(\ireg_m[12] ));
    NOR2 inf_abs1_a_2_I_15 (.A(sr_new[3]), .B(sr_new[4]), .Y(
        \DWACT_FINC_E_0[1] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I83_Y (.A(sum_17), .B(
        \un1_next_sum[17] ), .C(N520), .Y(N633));
    XA1B \sumreg_RNO[25]  (.A(N1055), .B(ADD_40x40_fast_I443_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[25] ));
    DFN1E1C0 \i_adj[11]  (.D(\inf_abs2_5[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[11]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I138_Y (.A(N614), .B(N611), .C(
        N610), .Y(N691));
    NOR3B \ireg_RNISRSK[9]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[9]_net_1 ), .Y(\un3_next_sum_m[9] ));
    DFN1E1C0 \ireg[11]  (.D(\next_ireg_3[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[11]_net_1 ));
    AND2 un1_sumreg_0_0_ADD_40x40_fast_I311_Y (.A(N798), .B(N814), .Y(
        N882));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I420_Y_0 (.A(sum_2_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I420_Y_0));
    DFN1C0 \state[3]  (.D(\state[6]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[3]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I158_Y (.A(I158_un1_Y), .B(N630), 
        .Y(N711));
    AO1 \ireg_RNI36EG1[14]  (.A(\ireg[14]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[14] ), .Y(
        \un1_next_sum_iv_1[14] ));
    MX2 \i_adj_RNO[17]  (.A(integral[23]), .B(\inf_abs2_a_0[17] ), .S(
        integral_1_0), .Y(\inf_abs2_5[17] ));
    DFN1E1C0 \i_adj[1]  (.D(\inf_abs2_5[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[1]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I80_Y (.A(N353), .B(N350), .C(
        N349), .Y(N388));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I86_Y (.A(N513_0), .B(N517), .C(
        N516), .Y(N636));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I236_Y (.A(I236_un1_Y), .B(N713), 
        .Y(N795));
    DFN1E1C0 \sumreg[3]  (.D(\next_sum[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_3));
    OR2 \state_RNIUSQN[4]  (.A(next_sum_1_sqmuxa_1), .B(
        next_sum_1_sqmuxa_2), .Y(\un1_next_sum_0_iv_0[25] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I358_un1_Y (.A(N794), .B(N810), 
        .C(N743), .Y(I358_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I220_Y (.A(N705), .B(N698), .C(
        N697), .Y(N779));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I256_Y (.A(I256_un1_Y), .B(N733), 
        .Y(N815));
    DFN1E1C0 \sumreg_1[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_1_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I382_Y_1 (.A(N762), .B(N777), .C(
        ADD_40x40_fast_I382_Y_0), .Y(ADD_40x40_fast_I382_Y_1));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I4_G0N (.A(\i_adj[4]_net_1 ), 
        .B(\i_adj[6]_net_1 ), .Y(N278));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I357_Y (.A(N791), .B(I304_un1_Y), 
        .C(I357_un1_Y), .Y(N1070));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I85_Y (.A(
        ADD_22x22_fast_I85_Y_0), .B(N354), .Y(N393));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I24_P0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[24] ), .C(\sumreg[24]_net_1 ), .Y(N544));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I142_Y (.A(N618), .B(N615), .C(
        N614), .Y(N695));
    DFN1C0 \state_0[1]  (.D(\state_RNIGTM6[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_0[1]_net_1 ));
    NOR3 inf_abs2_a_0_I_50 (.A(integral[22]), .B(integral[21]), .C(
        integral[23]), .Y(\DWACT_FINC_E[12] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I347_un1_Y_0 (.A(N698), .B(
        N690), .C(N788), .Y(ADD_40x40_fast_I347_un1_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I3_G0N (.A(\i_adj[5]_net_1 ), 
        .B(\i_adj[3]_net_1 ), .Y(N275));
    NOR3B \ireg_RNI9GKN[17]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[17]_net_1 ), .Y(\un3_next_sum_m[17] ));
    XNOR2 inf_abs1_a_2_I_9 (.A(sr_new[3]), .B(N_11_0), .Y(
        \inf_abs1_a_2[3] ));
    NOR3B inf_abs1_a_2_I_16 (.A(\DWACT_FINC_E_0[1] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[5]), .Y(N_8_0));
    NOR3B \ireg_RNION1B[7]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[7]_net_1 ), .C(integral_0_0), .Y(\ireg_m[7] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I355_un1_Y (.A(N872), .B(N819), 
        .Y(I355_un1_Y));
    AO1 next_ireg_3_0_ADD_22x22_fast_I46_Y (.A(N278), .B(N282), .C(
        N281), .Y(N351));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I13_G0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[15]_net_1 ), .Y(N305));
    AO1A \preg_RNIQRUV[12]  (.A(\preg[12]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[12] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I361_un1_Y (.A(N884), .B(
        \un1_next_sum[0] ), .Y(I361_un1_Y));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I350_un1_Y (.A(N809), .B(
        I318_un1_Y), .C(ADD_40x40_fast_I350_un1_Y_0), .Y(I350_un1_Y));
    VCC VCC_i (.Y(VCC));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I221_Y (.A(N698), .B(N706), .Y(
        N780));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I14_G0N (.A(
        \un1_next_sum_iv_1[14] ), .B(\un1_next_sum_iv_2[14] ), .C(
        sum_14), .Y(N513_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I116_Y (.A(N471), .B(I116_un1_Y), 
        .Y(N666));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I50_Y (.A(\sumreg[33]_net_1 ), 
        .B(\sumreg[32]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N600)
        );
    AND3 inf_abs1_a_2_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(
        \DWACT_FINC_E[4] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I6_G0N (.A(\un1_next_sum[6] ), 
        .B(sum_6), .Y(N489));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I309_Y (.A(N812), .B(N796), .Y(
        N880));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I418_Y (.A(N_228_1), .B(N_232), 
        .C(ADD_40x40_fast_I418_Y_0), .Y(\un1_sumreg[0] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I383_un1_Y (.A(
        ADD_40x40_fast_I383_un1_Y_0), .B(N848), .Y(I383_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I185_Y (.A(N661), .B(N657), .Y(
        N738));
    OA1 next_ireg_3_0_ADD_22x22_fast_I85_Y_0 (.A(\i_adj[4]_net_1 ), .B(
        \i_adj[2]_net_1 ), .C(N270), .Y(ADD_22x22_fast_I85_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I448_Y_0 (.A(
        \sumreg[30]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I448_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I107_Y (.A(N484), .B(N487), .Y(
        N657));
    AO1 next_ireg_3_0_ADD_22x22_fast_I129_Y_0 (.A(N384), .B(N377), .C(
        N376), .Y(ADD_22x22_fast_I129_Y_0));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I130_un1_Y (.A(N379), .B(N387), 
        .C(N394), .Y(I130_un1_Y));
    AO1 next_ireg_3_0_ADD_22x22_fast_I112_Y (.A(N387), .B(N394), .C(
        N386), .Y(N522));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I228_Y (.A(N713), .B(N706), .C(
        N705), .Y(N787));
    NOR3 inf_abs1_a_2_I_8 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2]), 
        .Y(N_11_0));
    XA1B \sumreg_RNO[26]  (.A(N1052), .B(ADD_40x40_fast_I444_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[26] ));
    AO1 \preg_RNI5I3J[7]  (.A(\preg[7]_net_1 ), .B(next_sum_1_sqmuxa_2)
        , .C(\ireg_m[7] ), .Y(\un1_next_sum_iv_1[7] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I454_Y_0 (.A(
        \sumreg[36]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I454_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I110_Y (.A(sum_2_d0), .B(
        \un1_next_sum[0] ), .C(N480), .Y(N660));
    XA1B \sumreg_RNO[17]  (.A(N1079), .B(ADD_40x40_fast_I435_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[17] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I286_un1_Y (.A(N707), .B(
        I230_un1_Y), .C(N774), .Y(I286_un1_Y));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I359_Y (.A(N795), .B(I308_un1_Y), 
        .C(I359_un1_Y), .Y(N1076));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I137_Y (.A(N613), .B(N609), .Y(
        N690));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I129_un1_Y_0 (.A(N377), .B(N385)
        , .Y(ADD_22x22_fast_I129_un1_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I453_Y_0 (.A(
        \sumreg[35]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I453_Y_0));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I48_Y (.A(\sumreg[33]_net_1 ), 
        .B(\sumreg[34]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N598)
        );
    NOR2A inf_abs1_a_2_I_25 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .Y(
        N_5));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I157_Y (.A(N629), .B(N633), .Y(
        N710));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I428_Y_0 (.A(
        \un1_next_sum_iv_1[10] ), .B(\un1_next_sum_iv_2[10] ), .C(
        sum_10), .Y(ADD_40x40_fast_I428_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I312_Y (.A(I312_un1_Y), .B(N799), 
        .Y(N883));
    DFN1E1C0 \preg[11]  (.D(\p_adj[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[11]_net_1 ));
    XA1B \sumreg_RNO[23]  (.A(N1061), .B(ADD_40x40_fast_I441_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[23] ));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I131_un1_Y (.A(N381), .B(N389), 
        .C(N396), .Y(I131_un1_Y));
    DFN1E1C0 \sumreg[22]  (.D(\next_sum[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_22));
    OR2 next_ireg_3_0_ADD_22x22_fast_I115_Y (.A(I115_un1_Y), .B(N392), 
        .Y(N531));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I5_P0N (.A(\un1_next_sum[5] ), 
        .B(sum_5), .Y(N487));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I66_un1_Y (.A(N543), .B(N547), 
        .Y(I66_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I20_G0N (.A(\un1_next_sum[20] )
        , .B(sum_20), .Y(N531_0));
    DFN1E1C0 \ireg[13]  (.D(\next_ireg_3[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[13]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I296_un1_Y (.A(N799), .B(N784), 
        .Y(I296_un1_Y));
    XA1B \sumreg_RNO[29]  (.A(N1043), .B(ADD_40x40_fast_I447_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[29] ));
    DFN1E1C0 \p_adj[8]  (.D(\inf_abs1_5[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[8]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I61_Y (.A(N334), .B(N330), .Y(
        N369));
    AX1D next_ireg_3_0_ADD_22x22_fast_I177_Y (.A(I124_un1_Y), .B(
        ADD_22x22_fast_I144_Y_2), .C(ADD_22x22_fast_I177_Y_0), .Y(
        \next_ireg_3[23] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I84_Y (.A(N357), .B(N354), .C(
        N353), .Y(N392));
    OR3 \preg_RNIQO7N1[18]  (.A(\un24_next_sum_m[18] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[18] ), .Y(
        \un1_next_sum_iv_2[18] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I240_Y (.A(I240_un1_Y), .B(N717), 
        .Y(N799));
    NOR3B \preg_RNIER18[8]  (.A(\state[5]_net_1 ), .B(\preg[8]_net_1 ), 
        .C(sr_new[12]), .Y(\preg_m[8] ));
    XNOR2 inf_abs1_a_2_I_7 (.A(sr_new[2]), .B(N_12), .Y(
        \inf_abs1_a_2[2] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I240_un1_Y (.A(N725), .B(N718), 
        .Y(I240_un1_Y));
    XNOR2 inf_abs2_a_0_I_17 (.A(integral[12]), .B(N_21), .Y(
        \inf_abs2_a_0[6] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_1_1 (.A(
        \i_adj[19]_net_1 ), .B(\i_adj[17]_net_1 ), .Y(N_14_1));
    NOR3B \ireg_RNIQPSK[7]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[7]_net_1 ), .Y(\un3_next_sum_m[7] ));
    DFN1E1C0 \sumreg[12]  (.D(\next_sum[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_12));
    DFN1E1C0 \ireg[15]  (.D(\next_ireg_3[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[15]_net_1 ));
    XA1B \sumreg_RNO[1]  (.A(N666), .B(ADD_40x40_fast_I419_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[1] ));
    AX1D next_ireg_3_0_ADD_22x22_fast_I179_Y (.A(N_12_0), .B(
        ADD_22x22_fast_I142_Y_0_1), .C(ADD_22x22_fast_I179_Y_0), .Y(
        \next_ireg_3[25] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I97_Y (.A(N499), .B(N502), .Y(
        N647));
    NOR2B \state_RNIGTM6[0]  (.A(sum_rdy), .B(sum_enable), .Y(
        \state_RNIGTM6[0]_net_1 ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I8_P0N (.A(\i_adj[10]_net_1 ), .B(
        \i_adj[8]_net_1 ), .Y(N291));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I280_un1_Y (.A(N694), .B(N686), 
        .C(N783), .Y(I280_un1_Y));
    DFN1E1C0 \sumreg_2[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIRSTG[6]_net_1 ), .Q(sum_2_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I7_P0N (.A(\i_adj[9]_net_1 ), .B(
        \i_adj[7]_net_1 ), .Y(N288));
    NOR3 inf_abs1_a_2_I_18 (.A(sr_new[3]), .B(sr_new[5]), .C(sr_new[4])
        , .Y(\DWACT_FINC_E_0[2] ));
    XNOR2 inf_abs1_a_2_I_26 (.A(sr_new[9]), .B(N_5), .Y(
        \inf_abs1_a_2[9] ));
    
endmodule


module sig_gen_1(
       vd_done,
       n_rst_c,
       clk_c,
       sig_old_i_0,
       sig_prev
    );
input  vd_done;
input  n_rst_c;
input  clk_c;
output sig_old_i_0;
output sig_prev;

    wire sig_prev_i, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(clk_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev_inst_1 (.D(vd_done), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(sig_prev));
    INV sig_old_RNO (.A(sig_prev), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module spi_stp_12s_1_3(
       cur_vd,
       N_29,
       din_33_c,
       n_rst_c,
       sck_12_c
    );
output [11:0] cur_vd;
input  N_29;
input  din_33_c;
input  n_rst_c;
input  sck_12_c;

    wire GND, VCC;
    
    DFN1E0C0 \sr[7]  (.D(cur_vd[6]), .CLK(sck_12_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[7]));
    DFN1E0C0 \sr[5]  (.D(cur_vd[4]), .CLK(sck_12_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[5]));
    DFN1E0C0 \sr[10]  (.D(cur_vd[9]), .CLK(sck_12_c), .CLR(n_rst_c), 
        .E(N_29), .Q(cur_vd[10]));
    DFN1E0C0 \sr[8]  (.D(cur_vd[7]), .CLK(sck_12_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[8]));
    DFN1E0C0 \sr[3]  (.D(cur_vd[2]), .CLK(sck_12_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[3]));
    DFN1E0C0 \sr[1]  (.D(cur_vd[0]), .CLK(sck_12_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[1]));
    DFN1E0C0 \sr[2]  (.D(cur_vd[1]), .CLK(sck_12_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[2]));
    DFN1E0C0 \sr[9]  (.D(cur_vd[8]), .CLK(sck_12_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[9]));
    VCC VCC_i (.Y(VCC));
    DFN1E0C0 \sr[11]  (.D(cur_vd[10]), .CLK(sck_12_c), .CLR(n_rst_c), 
        .E(N_29), .Q(cur_vd[11]));
    DFN1E0C0 \sr[0]  (.D(din_33_c), .CLK(sck_12_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[0]));
    GND GND_i (.Y(GND));
    DFN1E0C0 \sr[6]  (.D(cur_vd[5]), .CLK(sck_12_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[6]));
    DFN1E0C0 \sr[4]  (.D(cur_vd[3]), .CLK(sck_12_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[4]));
    
endmodule


module sig_gen_10_1(
       cs_i_1,
       n_rst_c,
       sck_12_c,
       vd_done
    );
input  cs_i_1;
input  n_rst_c;
input  sck_12_c;
output vd_done;

    wire sig_prev_i, sig_prev_net_1, sig_old_i_0, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(sck_12_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev (.D(cs_i_1), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        sig_prev_net_1));
    INV sig_old_RNO (.A(sig_prev_net_1), .Y(sig_prev_i));
    NOR2B sig_old_RNIALTK (.A(sig_prev_net_1), .B(sig_old_i_0), .Y(
        vd_done));
    GND GND_i (.Y(GND));
    
endmodule


module spi_ctl_12s_1(
       n_rst_c,
       sck_12_c,
       N_29,
       cs_i_1,
       cs_i_1_i
    );
input  n_rst_c;
input  sck_12_c;
output N_29;
output cs_i_1;
output cs_i_1_i;

    wire cnt_n6_i_o2_0, \cnt[5]_net_1 , \cnt[4]_net_1 , cnt_m1_0_a2_0, 
        \cnt[14]_net_1 , \cnt[13]_net_1 , cnt_m6_0_a2_6, cnt_m6_0_a2_0, 
        cnt_m5_0_a2_2, cnt_m6_0_a2_2, \cnt[7]_net_1 , \cnt[8]_net_1 , 
        \cnt[11]_net_1 , \cnt[10]_net_1 , cnt_m7_0_a2_4, cnt_m7_0_a2_3, 
        \cnt[6]_net_1 , cnt_m7_0_a2_1, \cnt[9]_net_1 , 
        state_tr0_0_a3_12, state_tr0_0_a3_6, state_tr0_0_a3_9, N_103, 
        state_tr0_0_a3_8, state_tr0_0_a3_4, state_tr0_0_a3_7, 
        state_tr0_0_a3_2, \cnt[0]_net_1 , \cnt[1]_net_1 , 
        state_tr0_0_a3_1, \cnt[15]_net_1 , \cnt[12]_net_1 , 
        vd_stp_en_i_a3_9, vd_stp_en_i_a3_4, vd_stp_en_i_a3_3, N_73, 
        vd_stp_en_i_a3_8, vd_stp_en_i_a3_2, vd_stp_en_i_a3_5, 
        cnt_m6_0_a2_5_6, cnt_m6_0_a2_5_0, cnt_m6_0_a2_5, 
        \cnt[2]_net_1 , cnt_m5_0_a2_3, cnt_m2_0_a2_0, \cnt[3]_net_1 , 
        cnt_m5_0_a2_1, cnt_m2_0_a2_2, cnt_m2_0_a2_1, N_74, 
        cnt_N_13_mux, N_34, N_32, cnt_N_7_mux_0_0, cnt_N_3_mux_0, 
        cnt_N_11_mux_2, cnt_N_15_mux, N_31, cnt_N_13_mux_0, N_30, 
        \state_RNO_2[0]_net_1 , N_26, N_24, N_22, N_20, N_18, N_96, 
        N_14, N_12, N_36, \cnt_RNO_3[6] , cnt_n10, d_N_3_mux_2, 
        \cnt_RNO_1_0[10] , cnt_n0, cnt_n15, cnt_n14, cnt_n13, N_72, 
        cnt_n12, cnt_n11, cnt_n9, N_38, GND, VCC;
    
    NOR2B \cnt_RNO_2[6]  (.A(\cnt[5]_net_1 ), .B(\cnt[4]_net_1 ), .Y(
        cnt_m2_0_a2_2));
    XA1A \cnt_RNO[8]  (.A(\cnt[8]_net_1 ), .B(N_36), .C(cs_i_1), .Y(
        N_12));
    NOR2B \cnt_RNO_3[10]  (.A(cnt_m5_0_a2_2), .B(cs_i_1), .Y(
        cnt_m7_0_a2_4));
    NOR3A \state_RNO_0[0]  (.A(state_tr0_0_a3_4), .B(\cnt[6]_net_1 ), 
        .C(\cnt[7]_net_1 ), .Y(state_tr0_0_a3_8));
    XA1A \cnt_RNO[2]  (.A(N_30), .B(\cnt[2]_net_1 ), .C(cs_i_1), .Y(
        N_24));
    DFN1C0 \cnt[2]  (.D(N_24), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[2]_net_1 ));
    DFN1C0 \cnt[8]  (.D(N_12), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[8]_net_1 ));
    DFN1C0 \cnt[1]  (.D(N_26), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[1]_net_1 ));
    DFN1C0 \cnt[11]  (.D(cnt_n11), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[11]_net_1 ));
    NOR3C \cnt_RNO_0[6]  (.A(cnt_m2_0_a2_1), .B(cnt_m2_0_a2_0), .C(
        cnt_m2_0_a2_2), .Y(cnt_N_7_mux_0_0));
    NOR3C \cnt_RNI1P4N2[2]  (.A(cnt_m5_0_a2_2), .B(cnt_m5_0_a2_1), .C(
        cnt_m5_0_a2_3), .Y(cnt_N_11_mux_2));
    NOR2B \cnt_RNO_1[15]  (.A(\cnt[14]_net_1 ), .B(\cnt[13]_net_1 ), 
        .Y(cnt_m1_0_a2_0));
    XA1A \cnt_RNO[3]  (.A(N_31), .B(\cnt[3]_net_1 ), .C(cs_i_1), .Y(
        N_22));
    OR2B \cnt_RNO_0[13]  (.A(cnt_N_13_mux), .B(\cnt[12]_net_1 ), .Y(
        N_72));
    NOR3B \state_RNO_6[0]  (.A(\cnt[5]_net_1 ), .B(N_103), .C(
        \cnt[4]_net_1 ), .Y(state_tr0_0_a3_9));
    NOR2B \cnt_RNIB9FL[11]  (.A(\cnt[11]_net_1 ), .B(\cnt[10]_net_1 ), 
        .Y(cnt_m6_0_a2_0));
    VCC VCC_i (.Y(VCC));
    OR2B \cnt_RNO_2[5]  (.A(\cnt[5]_net_1 ), .B(\cnt[4]_net_1 ), .Y(
        cnt_n6_i_o2_0));
    XA1 \cnt_RNO[1]  (.A(\cnt[0]_net_1 ), .B(\cnt[1]_net_1 ), .C(
        cs_i_1), .Y(N_26));
    DFN1C0 \cnt[6]  (.D(\cnt_RNO_3[6] ), .CLK(sck_12_c), .CLR(n_rst_c), 
        .Q(\cnt[6]_net_1 ));
    NOR3C \cnt_RNO_0[15]  (.A(cnt_m1_0_a2_0), .B(\cnt[12]_net_1 ), .C(
        cnt_N_13_mux), .Y(cnt_N_3_mux_0));
    NOR3A \state_RNO_1[0]  (.A(state_tr0_0_a3_2), .B(\cnt[0]_net_1 ), 
        .C(\cnt[1]_net_1 ), .Y(state_tr0_0_a3_7));
    NOR2B \cnt_RNI12B51[4]  (.A(\cnt[4]_net_1 ), .B(cnt_m2_0_a2_0), .Y(
        cnt_m5_0_a2_3));
    DFN1C0 \cnt[4]  (.D(N_20), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[4]_net_1 ));
    DFN1C0 \cnt[9]  (.D(cnt_n9), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[9]_net_1 ));
    NOR2A \cnt_RNO[0]  (.A(cs_i_1), .B(\cnt[0]_net_1 ), .Y(cnt_n0));
    OA1C \cnt_RNO_1[5]  (.A(\cnt[4]_net_1 ), .B(N_32), .C(
        \cnt[5]_net_1 ), .Y(N_96));
    OR3C \cnt_RNO_0[14]  (.A(\cnt[12]_net_1 ), .B(\cnt[13]_net_1 ), .C(
        cnt_N_13_mux), .Y(N_74));
    DFN1C0 \cnt[0]  (.D(cnt_n0), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[0]_net_1 ));
    XA1A \cnt_RNO[4]  (.A(\cnt[4]_net_1 ), .B(N_32), .C(cs_i_1), .Y(
        N_20));
    NOR2 \state_RNO_4[0]  (.A(\cnt[10]_net_1 ), .B(\cnt[8]_net_1 ), .Y(
        state_tr0_0_a3_2));
    OR2B \cnt_RNIS9J33[7]  (.A(cnt_N_11_mux_2), .B(\cnt[7]_net_1 ), .Y(
        N_36));
    NOR2 \cnt_RNIM1TO[6]  (.A(\cnt[8]_net_1 ), .B(\cnt[6]_net_1 ), .Y(
        vd_stp_en_i_a3_3));
    DFN1C0 \state[0]  (.D(\state_RNO_2[0]_net_1 ), .CLK(sck_12_c), 
        .CLR(n_rst_c), .Q(cs_i_1));
    XA1 \cnt_RNO[6]  (.A(cnt_N_7_mux_0_0), .B(\cnt[6]_net_1 ), .C(
        cs_i_1), .Y(\cnt_RNO_3[6] ));
    XA1 \cnt_RNO[15]  (.A(\cnt[15]_net_1 ), .B(cnt_N_3_mux_0), .C(
        cs_i_1), .Y(cnt_n15));
    XA1A \cnt_RNO[9]  (.A(\cnt[9]_net_1 ), .B(N_38), .C(cs_i_1), .Y(
        cnt_n9));
    GND GND_i (.Y(GND));
    NOR2B \cnt_RNO_5[10]  (.A(\cnt[8]_net_1 ), .B(\cnt[9]_net_1 ), .Y(
        cnt_m7_0_a2_1));
    NOR2B \cnt_RNIGRSO[2]  (.A(\cnt[2]_net_1 ), .B(\cnt[6]_net_1 ), .Y(
        cnt_m5_0_a2_1));
    NOR3C \cnt_RNIE5QH1[9]  (.A(\cnt[9]_net_1 ), .B(\cnt[6]_net_1 ), 
        .C(cnt_m6_0_a2_2), .Y(cnt_m6_0_a2_5));
    DFN1C0 \cnt[13]  (.D(cnt_n13), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[13]_net_1 ));
    NOR3A \state_RNO_5[0]  (.A(state_tr0_0_a3_1), .B(\cnt[14]_net_1 ), 
        .C(\cnt[15]_net_1 ), .Y(state_tr0_0_a3_6));
    OR2A \cnt_RNO_0[9]  (.A(\cnt[8]_net_1 ), .B(N_36), .Y(N_38));
    DFN1C0 \cnt[7]  (.D(N_14), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[7]_net_1 ));
    NOR3C \state_RNO_2[0]  (.A(state_tr0_0_a3_6), .B(cs_i_1), .C(
        state_tr0_0_a3_9), .Y(state_tr0_0_a3_12));
    OR2A \cnt_RNI56B51[4]  (.A(\cnt[4]_net_1 ), .B(N_103), .Y(N_73));
    NOR3C \cnt_RNI6NSC2[10]  (.A(vd_stp_en_i_a3_2), .B(
        state_tr0_0_a3_1), .C(vd_stp_en_i_a3_5), .Y(vd_stp_en_i_a3_8));
    DFN1C0 \cnt[10]  (.D(cnt_n10), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[10]_net_1 ));
    NOR2 \cnt_RNICAFL[10]  (.A(\cnt[10]_net_1 ), .B(\cnt[12]_net_1 ), 
        .Y(vd_stp_en_i_a3_2));
    NOR2B \cnt_RNI9KSO_0[1]  (.A(\cnt[1]_net_1 ), .B(\cnt[0]_net_1 ), 
        .Y(cnt_m2_0_a2_0));
    NOR3C \cnt_RNO_1[11]  (.A(cnt_m6_0_a2_5_0), .B(\cnt[4]_net_1 ), .C(
        cnt_m5_0_a2_2), .Y(cnt_m6_0_a2_5_6));
    NOR3B \cnt_RNO[5]  (.A(N_34), .B(cs_i_1), .C(N_96), .Y(N_18));
    NOR3C \cnt_RNIJIQQ1[4]  (.A(cnt_m6_0_a2_0), .B(\cnt[4]_net_1 ), .C(
        cnt_m5_0_a2_2), .Y(cnt_m6_0_a2_6));
    NOR3 \cnt_RNIC0U11[15]  (.A(\cnt[14]_net_1 ), .B(\cnt[15]_net_1 ), 
        .C(\cnt[5]_net_1 ), .Y(vd_stp_en_i_a3_5));
    INV \state_RNIGSV6[0]  (.A(cs_i_1), .Y(cs_i_1_i));
    DFN1C0 \cnt[3]  (.D(N_22), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[3]_net_1 ));
    NOR2B \cnt_RNO_2[11]  (.A(\cnt[10]_net_1 ), .B(\cnt[2]_net_1 ), .Y(
        cnt_m6_0_a2_5_0));
    XA1A \cnt_RNO[14]  (.A(\cnt[14]_net_1 ), .B(N_74), .C(cs_i_1), .Y(
        cnt_n14));
    NOR2 \cnt_RNIO3TO[9]  (.A(\cnt[9]_net_1 ), .B(\cnt[7]_net_1 ), .Y(
        vd_stp_en_i_a3_4));
    NOR2B \cnt_RNIN2TO[7]  (.A(\cnt[7]_net_1 ), .B(\cnt[8]_net_1 ), .Y(
        cnt_m6_0_a2_2));
    OR2A \cnt_RNIMCPH1[3]  (.A(\cnt[3]_net_1 ), .B(N_31), .Y(N_32));
    OR2B \cnt_RNI9KSO[1]  (.A(\cnt[1]_net_1 ), .B(\cnt[0]_net_1 ), .Y(
        N_30));
    NOR3C \cnt_RNIJB5N2[4]  (.A(vd_stp_en_i_a3_4), .B(vd_stp_en_i_a3_3)
        , .C(N_73), .Y(vd_stp_en_i_a3_9));
    XNOR2 \cnt_RNO_1[10]  (.A(\cnt[10]_net_1 ), .B(\cnt[4]_net_1 ), .Y(
        \cnt_RNO_1_0[10] ));
    NOR3C \cnt_RNO_4[10]  (.A(\cnt[7]_net_1 ), .B(\cnt[6]_net_1 ), .C(
        cnt_m7_0_a2_1), .Y(cnt_m7_0_a2_3));
    NOR3B \cnt_RNO_0[11]  (.A(cnt_m6_0_a2_5), .B(cnt_m6_0_a2_5_6), .C(
        N_30), .Y(cnt_N_13_mux_0));
    XA1 \cnt_RNO[11]  (.A(\cnt[11]_net_1 ), .B(cnt_N_13_mux_0), .C(
        cs_i_1), .Y(cnt_n11));
    NOR3B \cnt_RNI0OVH4[4]  (.A(cnt_m6_0_a2_6), .B(cnt_m6_0_a2_5), .C(
        N_31), .Y(cnt_N_13_mux));
    NOR3B \cnt_RNO_2[10]  (.A(cnt_m7_0_a2_4), .B(cnt_m7_0_a2_3), .C(
        N_31), .Y(cnt_N_15_mux));
    NOR2 \cnt_RNIECFL[11]  (.A(\cnt[11]_net_1 ), .B(\cnt[13]_net_1 ), 
        .Y(state_tr0_0_a3_1));
    OR3C \state_RNO[0]  (.A(state_tr0_0_a3_8), .B(state_tr0_0_a3_7), 
        .C(state_tr0_0_a3_12), .Y(\state_RNO_2[0]_net_1 ));
    MX2B \cnt_RNO[10]  (.A(d_N_3_mux_2), .B(\cnt_RNO_1_0[10] ), .S(
        cnt_N_15_mux), .Y(cnt_n10));
    DFN1C0 \cnt[15]  (.D(cnt_n15), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[15]_net_1 ));
    OR2 \cnt_RNO_0[5]  (.A(cnt_n6_i_o2_0), .B(N_32), .Y(N_34));
    OR2A \cnt_RNIVVA51[2]  (.A(\cnt[2]_net_1 ), .B(N_30), .Y(N_31));
    AO1B \state_RNI9V1B5[0]  (.A(vd_stp_en_i_a3_9), .B(
        vd_stp_en_i_a3_8), .C(cs_i_1), .Y(N_29));
    NOR2B \cnt_RNO_1[6]  (.A(\cnt[2]_net_1 ), .B(\cnt[3]_net_1 ), .Y(
        cnt_m2_0_a2_1));
    NOR2B \cnt_RNIGRSO[3]  (.A(\cnt[3]_net_1 ), .B(\cnt[5]_net_1 ), .Y(
        cnt_m5_0_a2_2));
    NOR2B \cnt_RNO_0[10]  (.A(\cnt[10]_net_1 ), .B(cs_i_1), .Y(
        d_N_3_mux_2));
    NOR2 \state_RNO_3[0]  (.A(\cnt[9]_net_1 ), .B(\cnt[12]_net_1 ), .Y(
        state_tr0_0_a3_4));
    DFN1C0 \cnt[5]  (.D(N_18), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[5]_net_1 ));
    XA1A \cnt_RNO[13]  (.A(\cnt[13]_net_1 ), .B(N_72), .C(cs_i_1), .Y(
        cnt_n13));
    NOR2 \cnt_RNIDOSO[3]  (.A(\cnt[3]_net_1 ), .B(\cnt[2]_net_1 ), .Y(
        N_103));
    XA1 \cnt_RNO[12]  (.A(\cnt[12]_net_1 ), .B(cnt_N_13_mux), .C(
        cs_i_1), .Y(cnt_n12));
    DFN1C0 \cnt[12]  (.D(cnt_n12), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[12]_net_1 ));
    XA1 \cnt_RNO[7]  (.A(\cnt[7]_net_1 ), .B(cnt_N_11_mux_2), .C(
        cs_i_1), .Y(N_14));
    DFN1C0 \cnt[14]  (.D(cnt_n14), .CLK(sck_12_c), .CLR(n_rst_c), .Q(
        \cnt[14]_net_1 ));
    
endmodule


module spi_rx_12s_1(
       cur_vd,
       vd_done,
       cs_i_1_i,
       sck_12_c,
       n_rst_c,
       din_33_c
    );
output [11:0] cur_vd;
output vd_done;
output cs_i_1_i;
input  sck_12_c;
input  n_rst_c;
input  din_33_c;

    wire N_29, cs_i_1, GND, VCC;
    
    spi_stp_12s_1_3 VD_STP (.cur_vd({cur_vd[11], cur_vd[10], cur_vd[9], 
        cur_vd[8], cur_vd[7], cur_vd[6], cur_vd[5], cur_vd[4], 
        cur_vd[3], cur_vd[2], cur_vd[1], cur_vd[0]}), .N_29(N_29), 
        .din_33_c(din_33_c), .n_rst_c(n_rst_c), .sck_12_c(sck_12_c));
    sig_gen_10_1 SPI_RDYSIG (.cs_i_1(cs_i_1), .n_rst_c(n_rst_c), 
        .sck_12_c(sck_12_c), .vd_done(vd_done));
    VCC VCC_i (.Y(VCC));
    spi_ctl_12s_1 SPICTL (.n_rst_c(n_rst_c), .sck_12_c(sck_12_c), 
        .N_29(N_29), .cs_i_1(cs_i_1), .cs_i_1_i(cs_i_1_i));
    GND GND_i (.Y(GND));
    
endmodule


module integral_calc_13s_0_4_0(
       sr_new,
       sr_old,
       sr_new_1_0,
       sr_new_0_0,
       integral,
       integral_i,
       integral_0_0,
       integral_1_0,
       calc_int,
       N_46_1,
       n_rst_c,
       clk_c
    );
input  [12:0] sr_new;
input  [12:0] sr_old;
input  sr_new_1_0;
input  sr_new_0_0;
output [25:6] integral;
output [25:24] integral_i;
output integral_0_0;
output integral_1_0;
input  calc_int;
output N_46_1;
input  n_rst_c;
input  clk_c;

    wire \un1_integ[25] , \un1_next_int_0_iv_0[13] , next_int_1_sqmuxa, 
        next_int_0_sqmuxa_1, N_46_1_0, \state[1]_net_1 , 
        \state[0]_net_1 , N_12, N_10, \DWACT_FINC_E[0] , N_5, 
        \DWACT_FINC_E[4] , N_2, \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , 
        N_12_0, N_10_0, \DWACT_FINC_E_0[0] , N_5_0, 
        \DWACT_FINC_E_0[4] , N_2_0, \DWACT_FINC_E_0[7] , 
        \DWACT_FINC_E_0[6] , ADD_26x26_fast_I255_Y_0, 
        \un1_next_int_0_iv[13] , ADD_26x26_fast_I254_Y_0, 
        ADD_26x26_fast_I253_Y_0, ADD_26x26_fast_I252_Y_0, 
        ADD_26x26_fast_I249_Y_0, ADD_26x26_fast_I247_Y_0, 
        ADD_26x26_fast_I204_Y_3, N517, N502, ADD_26x26_fast_I204_Y_2, 
        N455, N448, ADD_26x26_fast_I204_Y_1, ADD_26x26_fast_I204_Y_0, 
        N398, ADD_26x26_fast_I205_Y_3, N504, N519, 
        ADD_26x26_fast_I205_Y_2, N450, N457, ADD_26x26_fast_I205_Y_1, 
        N397, N400, ADD_26x26_fast_I205_Y_0, ADD_26x26_fast_I248_Y_0, 
        ADD_26x26_fast_I250_Y_0, ADD_26x26_fast_I251_Y_0, 
        ADD_26x26_fast_I206_Y_2, ADD_26x26_fast_I206_un1_Y_0, N522, 
        ADD_26x26_fast_I206_Y_1, N459, N452, ADD_26x26_fast_I206_Y_0, 
        N402, N399, ADD_26x26_fast_I245_Y_0, ADD_26x26_fast_I207_Y_2, 
        ADD_26x26_fast_I207_un1_Y_0, N524, ADD_26x26_fast_I207_Y_1, 
        N454, N461, ADD_26x26_fast_I207_Y_0, N401, N404, 
        ADD_26x26_fast_I210_Y_1, N529, N514, ADD_26x26_fast_I210_Y_0, 
        N467, N460, ADD_26x26_fast_I212_Y_0, N533, N518, 
        ADD_26x26_fast_I242_Y_0, \un2_next_int_m[12] , 
        \un1_next_int_iv_0[12] , ADD_26x26_fast_I244_Y_0, 
        ADD_26x26_fast_I243_Y_0, ADD_26x26_fast_I211_Y_0, N462, N469, 
        ADD_26x26_fast_I208_Y_1, ADD_26x26_fast_I208_un1_Y_0, N526, 
        ADD_26x26_fast_I208_Y_0, N463, N456, ADD_26x26_fast_I209_Y_1, 
        ADD_26x26_fast_I209_un1_Y_0, N528, ADD_26x26_fast_I209_Y_0, 
        N458, N465, ADD_26x26_fast_I204_un1_Y_0, 
        ADD_26x26_fast_I239_Y_0, \un2_next_int_m[9] , 
        \un1_next_int_iv_1[9] , ADD_26x26_fast_I240_Y_0, 
        \un1_next_int[10] , ADD_26x26_fast_I211_Y_1_0, N470, 
        ADD_26x26_fast_I213_un1_Y_0, N482, N490, 
        \state_RNICBRB4[0]_net_1 , N483, I160_un1_Y, N506, N487, 
        I162_un1_Y, N510, N485, I161_un1_Y, N508, N543, N512, 
        ADD_26x26_fast_I237_Y_0, \un2_next_int_m[7] , 
        \un1_next_int_iv_1[7] , ADD_26x26_fast_I236_Y_0, 
        \un1_next_int[6] , ADD_26x26_fast_I235_Y_0, \integ[5]_net_1 , 
        \un1_next_int[5] , ADD_26x26_fast_I233_Y_0, \integ[3]_net_1 , 
        \un1_next_int[3] , ADD_26x26_fast_I77_Y_0, 
        \un1_next_int_iv_0[11] , \inf_abs1[11]_net_1 , 
        \un1_next_int_iv_0[10] , \inf_abs1[10]_net_1 , 
        \un1_next_int_iv_0[8] , \inf_abs1[8]_net_1 , 
        \un1_next_int_iv_0[4] , \inf_abs1[4]_net_1 , 
        \un1_next_int_iv_0[6] , \inf_abs1[6]_net_1 , 
        ADD_26x26_fast_I230_Y_0, \integ[0]_net_1 , N_3, 
        \inf_abs0_m[9] , \un18_next_int_m[9] , \inf_abs1_m[9] , 
        \inf_abs1_a_1[12] , \un1_next_int_iv_1[0] , \inf_abs1_m[0] , 
        \un18_next_int_m[0] , \inf_abs0_m[0] , \inf_abs0_m[7] , 
        \un18_next_int_m[7] , \inf_abs1_m[7] , \un1_next_int_iv_1[5] , 
        \inf_abs0_m[5] , \un18_next_int_m[5] , \inf_abs1_m[5] , 
        \un1_next_int_iv_0[2] , \inf_abs1[2]_net_1 , 
        \un1_next_int_iv_1[3] , \inf_abs1_m[3] , \un18_next_int_m[3] , 
        \inf_abs0_m[3] , \un1_next_int_iv_1[1] , 
        \un1_next_int_iv_0[1] , \inf_abs0_m[1] , \inf_abs1[1]_net_1 , 
        ADD_26x26_fast_I211_Y_1, ADD_26x26_fast_I211_un1_Y_0, N531, 
        \un2_next_int_m[3] , \un2_next_int_m[5] , \inf_abs0_m[10] , 
        \un2_next_int_m[10] , \un1_next_int[1] , \un2_next_int_m[1] , 
        \un2_next_int_m[0] , \un1_next_int[2] , \inf_abs0_m[2] , 
        \un2_next_int_m[2] , \un1_next_int[4] , \inf_abs0_m[4] , 
        \un2_next_int_m[4] , \inf_abs0_m[6] , \un2_next_int_m[6] , 
        \un1_next_int[8] , \inf_abs0_m[8] , \un2_next_int_m[8] , 
        \state_RNIKDT9C[0]_net_1 , \inf_abs0_m[11] , 
        \un2_next_int_m[11] , \un1_integ[9] , I194_un1_Y, 
        \un1_integ[14] , N523, I189_un1_Y, I212_un1_Y, N534, N442, 
        I213_un1_Y, N520, N635, I186_un1_Y, \un1_integ[21] , 
        I176_un1_Y, \un1_integ[13] , N525, I190_un1_Y, \un1_integ[17] , 
        \un1_integ[16] , \un1_integ[20] , I178_un1_Y, \un1_integ[6] , 
        \un1_integ[15] , N521, I188_un1_Y, \un1_integ[12] , N527, 
        I191_un1_Y, \un1_integ[1] , \integ[1]_net_1 , \un1_integ[5] , 
        \un1_integ[0] , I204_un1_Y, \un1_integ[24] , I205_un1_Y, 
        \un1_integ[3] , N491, \un1_integ[7] , \un1_integ[18] , 
        \un1_integ[19] , I210_un1_Y, \un1_integ[23] , I172_un1_Y, 
        \un1_integ[2] , \integ[2]_net_1 , N493, \un1_integ[10] , 
        I193_un1_Y, \un1_integ[22] , I174_un1_Y, \un1_integ[11] , N649, 
        \un1_integ[8] , N658, \un1_integ[4] , \integ[4]_net_1 , N530, 
        N478, N486, N481, I158_un1_Y, I195_un1_Y, I150_un1_Y, N473, 
        N474, N466, N468, \state_RNO_1[0] , \state_RNO_2[1] , 
        I144_un1_Y, N475, N408, N409, N412, I146_un1_Y, N477, N436, 
        I118_un1_Y, I163_un1_Y, N426, N338, N427, N339, N431, N333, 
        N336, N488, N439, N435, N327, N421, N425, N345, N429, N323, 
        N326, N440, N437, N324, N441, N433, I110_un1_Y, N428, 
        I60_un1_Y, N432, N430, N332, N438, N434, I120_un1_Y, N476, 
        N403, N329, N350, N351, N424, N341, N344, I64_un1_Y, 
        I106_un1_Y, \inf_abs0[4]_net_1 , \inf_abs0[6]_net_1 , 
        \inf_abs0[8]_net_1 , \inf_abs0[11]_net_1 , \inf_abs0_a_0[4] , 
        \inf_abs0_a_0[6] , \inf_abs0_a_0[8] , \inf_abs0_a_0[11] , 
        \inf_abs1_a_1[4] , \inf_abs1_a_1[6] , \inf_abs1_a_1[8] , 
        \inf_abs1_a_1[11] , \inf_abs0[2]_net_1 , \inf_abs0_a_0[2] , 
        \inf_abs1_a_1[1] , \inf_abs1_a_1[2] , \inf_abs0_a_0[1] , N317, 
        N321, N320, N318, N416, N413, N410, N406, N353, N417, N354, 
        N464, N411, N415, N419, N414, N471, N422, N418, I104_un1_Y, 
        N423, N480, N479, I148_un1_Y, \inf_abs1_a_1[10] , 
        \inf_abs0[10]_net_1 , \inf_abs0_a_0[10] , N348, N347, N484, 
        N420, N405, N407, \inf_abs0_a_0[12] , \inf_abs0_a_0[5] , 
        \inf_abs1_a_1[5] , \inf_abs1_a_1[9] , \inf_abs0_a_0[9] , 
        \inf_abs1_a_1[7] , \inf_abs0_a_0[7] , \inf_abs1_a_1[3] , 
        \inf_abs0_a_0[3] , N_3_0, \DWACT_FINC_E[2] , \DWACT_FINC_E[5] , 
        N_4, \DWACT_FINC_E[3] , N_6, N_7, N_8, \DWACT_FINC_E[1] , N_9, 
        N_11, N_3_1, \DWACT_FINC_E_0[2] , \DWACT_FINC_E_0[5] , N_4_0, 
        \DWACT_FINC_E_0[3] , N_6_0, N_7_0, N_8_0, \DWACT_FINC_E_0[1] , 
        N_9_0, N_11_0, GND, VCC;
    
    AO1 un1_integ_0_0_ADD_26x26_fast_I56_Y (.A(N341), .B(N345), .C(
        N344), .Y(N424));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I148_un1_Y (.A(N419), .B(N423), 
        .C(N479), .Y(I148_un1_Y));
    NOR2 inf_abs1_a_1_I_15 (.A(sr_old[3]), .B(sr_old[4]), .Y(
        \DWACT_FINC_E[1] ));
    XNOR2 inf_abs1_a_1_I_23 (.A(sr_old[8]), .B(N_6), .Y(
        \inf_abs1_a_1[8] ));
    DFN1C0 \state[0]  (.D(\state_RNO_1[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[0]_net_1 ));
    XNOR2 inf_abs1_a_1_I_17 (.A(sr_old[6]), .B(N_8), .Y(
        \inf_abs1_a_1[6] ));
    DFN1E0C0 \integ[13]  (.D(\un1_integ[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[13]));
    DFN1E0C0 \integ[24]  (.D(\un1_integ[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[24]));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I245_Y_0 (.A(integral[15]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I245_Y_0));
    OA1A \state_RNIO4IK5[1]  (.A(sr_old[12]), .B(\inf_abs1_a_1[12] ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[12] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I61_Y (.A(N336), .B(N339), .Y(
        N429));
    NOR2B \state_RNILCQR1[0]  (.A(\inf_abs0[2]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[2] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I7_P0N (.A(\un2_next_int_m[7] ), 
        .B(\un1_next_int_iv_1[7] ), .C(integral[7]), .Y(N339));
    XA1A \state_RNIAG5D3[1]  (.A(sr_old[12]), .B(\inf_abs1[4]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[4] ));
    NOR3B inf_abs0_a_0_I_19 (.A(\DWACT_FINC_E_0[2] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[6]), .Y(N_7_0));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I248_Y_0 (.A(integral[18]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I248_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I172_un1_Y (.A(N506), .B(N521), 
        .Y(I172_un1_Y));
    NOR3B inf_abs0_a_0_I_16 (.A(\DWACT_FINC_E_0[1] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[5]), .Y(N_8_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I41_Y (.A(integral[16]), .B(
        integral[17]), .C(\un1_next_int_0_iv_0[13] ), .Y(N409));
    OA1 un1_integ_0_0_ADD_26x26_fast_I204_un1_Y (.A(N533), .B(
        I194_un1_Y), .C(ADD_26x26_fast_I204_un1_Y_0), .Y(I204_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I86_Y (.A(N404), .B(N408), .Y(
        N457));
    NOR3B \state_RNIOAH03[0]  (.A(sr_new_1_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[9] ), .Y(\un2_next_int_m[9] ));
    OR2 \state_RNISBO51_0[1]  (.A(next_int_1_sqmuxa), .B(
        next_int_0_sqmuxa_1), .Y(\un1_next_int_0_iv[13] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I98_Y (.A(N420), .B(N417), .C(
        N416), .Y(N469));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I176_un1_Y (.A(N525), .B(N510), 
        .Y(I176_un1_Y));
    OA1 un1_integ_0_0_ADD_26x26_fast_I158_un1_Y (.A(N436), .B(
        I118_un1_Y), .C(N482), .Y(I158_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I150_un1_Y (.A(N481), .B(N474), 
        .Y(I150_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I51_Y (.A(N354), .B(N351), .Y(
        N419));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y (.A(
        ADD_26x26_fast_I230_Y_0), .B(\state_RNICBRB4[0]_net_1 ), .Y(
        \un1_integ[0] ));
    NOR2B inf_abs1_a_1_I_34 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .Y(N_2_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I144_un1_Y (.A(N475), .B(N468), 
        .Y(I144_un1_Y));
    NOR3A \state_RNI08441[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .C(sr_old[3]), .Y(\un18_next_int_m[3] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I253_Y (.A(I172_un1_Y), .B(
        ADD_26x26_fast_I206_Y_2), .C(ADD_26x26_fast_I253_Y_0), .Y(
        \un1_integ[23] ));
    NOR2B \state_RNIHMBM[0]  (.A(sr_new[7]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[7] ));
    DFN1E0C0 \integ[21]  (.D(\un1_integ[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[21]));
    XNOR2 inf_abs1_a_1_I_7 (.A(sr_old[2]), .B(N_12_0), .Y(
        \inf_abs1_a_1[2] ));
    DFN1E0C0 \integ_1[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral_1_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I190_un1_Y (.A(N487), .B(
        I162_un1_Y), .C(N526), .Y(I190_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I146_Y (.A(I146_un1_Y), .B(N469), 
        .Y(N523));
    AO1 un1_integ_0_0_ADD_26x26_fast_I142_Y (.A(N466), .B(N473), .C(
        N465), .Y(N519));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I244_Y_0 (.A(integral[14]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I244_Y_0));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I231_Y (.A(\un1_next_int[1] ), 
        .B(\integ[1]_net_1 ), .C(N442), .Y(\un1_integ[1] ));
    AND3 inf_abs1_a_1_I_24 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E_0[4] ));
    OR2 \state_RNISS287[0]  (.A(\un1_next_int_iv_1[5] ), .B(
        \un2_next_int_m[5] ), .Y(\un1_next_int[5] ));
    XNOR2 inf_abs1_a_1_I_32 (.A(sr_old[11]), .B(N_3_0), .Y(
        \inf_abs1_a_1[11] ));
    OR2 \state_RNI3J5U2[1]  (.A(\un1_next_int_iv_0[1] ), .B(
        \inf_abs0_m[1] ), .Y(\un1_next_int_iv_1[1] ));
    DFN1E0C0 \integ[15]  (.D(\un1_integ[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[15]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I213_un1_Y (.A(
        ADD_26x26_fast_I213_un1_Y_0), .B(N520), .Y(I213_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I103_Y (.A(N421), .B(N425), .Y(
        N474));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I125_Y (.A(N456), .B(N448), .Y(
        N502));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_1 (.A(
        ADD_26x26_fast_I209_un1_Y_0), .B(N528), .C(
        ADD_26x26_fast_I209_Y_0), .Y(ADD_26x26_fast_I209_Y_1));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I97_Y (.A(N415), .B(N419), .Y(
        N468));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I77_Y (.A(
        ADD_26x26_fast_I77_Y_0), .B(N399), .Y(N448));
    AO1 un1_integ_0_0_ADD_26x26_fast_I94_Y (.A(N416), .B(N413), .C(
        N412), .Y(N465));
    XA1A \state_RNITG8K2[1]  (.A(sr_old[12]), .B(\inf_abs1[2]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[2] ));
    NOR2 inf_abs0_a_0_I_6 (.A(sr_new[0]), .B(sr_new[1]), .Y(N_12));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I81_Y (.A(N399), .B(N403), .Y(
        N452));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I151_Y (.A(N482), .B(N474), .Y(
        N528));
    AND3 inf_abs1_a_1_I_22 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_6));
    AO1 un1_integ_0_0_ADD_26x26_fast_I74_Y (.A(N318), .B(
        \state_RNICBRB4[0]_net_1 ), .C(N317), .Y(N442));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I238_Y (.A(\un1_next_int[8] ), 
        .B(integral[8]), .C(N658), .Y(\un1_integ[8] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I121_Y (.A(N441), .B(
        \state_RNICBRB4[0]_net_1 ), .C(N440), .Y(N493));
    NOR3 inf_abs0_a_0_I_10 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2])
        , .Y(\DWACT_FINC_E[0] ));
    XA1A \state_RNIN3IK5[1]  (.A(sr_old[12]), .B(\inf_abs1[10]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[10] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I5_P0N (.A(\integ[5]_net_1 ), .B(
        \un1_next_int[5] ), .Y(N333));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I236_Y_0 (.A(integral[6]), .B(
        \un1_next_int[6] ), .Y(ADD_26x26_fast_I236_Y_0));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I246_Y (.A(
        \un1_next_int_0_iv_0[13] ), .B(integral[16]), .C(N635), .Y(
        \un1_integ[16] ));
    NOR2B \state_RNIBGBM[0]  (.A(sr_new[1]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[1] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I252_Y_0 (.A(integral[22]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I252_Y_0));
    MX2 \inf_abs0[6]  (.A(sr_new[6]), .B(\inf_abs0_a_0[6] ), .S(
        sr_new_0_0), .Y(\inf_abs0[6]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I39_Y (.A(integral[17]), .B(
        integral[18]), .C(\un1_next_int_0_iv_0[13] ), .Y(N407));
    OA1B un1_integ_0_0_ADD_26x26_fast_I32_Y (.A(integral[21]), .B(
        integral[20]), .C(\un1_next_int_0_iv_0[13] ), .Y(N400));
    OR3 un1_integ_0_0_ADD_26x26_fast_I213_Y (.A(I186_un1_Y), .B(N519), 
        .C(I213_un1_Y), .Y(N635));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I194_un1_Y (.A(N534), .B(N442), 
        .Y(I194_un1_Y));
    NOR2A inf_abs0_a_0_I_11 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .Y(
        N_10));
    OR3 \state_RNI7AOSB[0]  (.A(\inf_abs0_m[10] ), .B(
        \un1_next_int_iv_0[10] ), .C(\un2_next_int_m[10] ), .Y(
        \un1_next_int[10] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I211_Y_1_0 (.A(N462), .B(N470), 
        .Y(ADD_26x26_fast_I211_Y_1_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I100_Y (.A(N422), .B(N419), .C(
        N418), .Y(N471));
    OR3 un1_integ_0_0_ADD_26x26_fast_I12_P0N (.A(\un2_next_int_m[12] ), 
        .B(\un1_next_int_iv_0[12] ), .C(integral[12]), .Y(N354));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I10_G0N (.A(integral[10]), .B(
        \un1_next_int[10] ), .Y(N347));
    NOR2B \state_RNISM6K4[1]  (.A(\inf_abs1_a_1[9] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[9] ));
    DFN1E0C0 \integ[12]  (.D(\un1_integ[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[12]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I109_Y (.A(N427), .B(N431), .Y(
        N480));
    XNOR2 inf_abs1_a_1_I_35 (.A(sr_old[12]), .B(N_2_0), .Y(
        \inf_abs1_a_1[12] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I205_Y_0 (.A(integral[22]), .B(
        integral[23]), .C(\un1_next_int_0_iv[13] ), .Y(
        ADD_26x26_fast_I205_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I115_Y (.A(N433), .B(N437), .Y(
        N486));
    OA1 un1_integ_0_0_ADD_26x26_fast_I12_G0N (.A(\un2_next_int_m[12] ), 
        .B(\un1_next_int_iv_0[12] ), .C(integral[12]), .Y(N353));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_0 (.A(N463), .B(N456), .C(
        N455), .Y(ADD_26x26_fast_I208_Y_0));
    NOR2 \state_RNIB7PP[0]  (.A(\state[1]_net_1 ), .B(\state[0]_net_1 )
        , .Y(N_46_1));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I111_Y (.A(N433), .B(N429), .Y(
        N482));
    NOR2A inf_abs1_a_1_I_25 (.A(\DWACT_FINC_E_0[4] ), .B(sr_old[8]), 
        .Y(N_5_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I2_P0N (.A(\integ[2]_net_1 ), .B(
        \un1_next_int[2] ), .Y(N324));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I250_Y_0 (.A(integral[20]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I250_Y_0));
    NOR3A inf_abs1_a_1_I_27 (.A(\DWACT_FINC_E_0[4] ), .B(sr_old[8]), 
        .C(sr_old[9]), .Y(N_4));
    DFN1E0C0 \integ[10]  (.D(\un1_integ[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[10]));
    OA1 un1_integ_0_0_ADD_26x26_fast_I188_un1_Y (.A(N483), .B(
        I160_un1_Y), .C(N522), .Y(I188_un1_Y));
    NOR3B \state_RNILI6B2[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[5] ), .Y(\un2_next_int_m[5] ));
    MX2 \inf_abs1[10]  (.A(sr_old[10]), .B(\inf_abs1_a_1[10] ), .S(
        sr_old[12]), .Y(\inf_abs1[10]_net_1 ));
    NOR3A \state_RNIT4441_0[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .C(sr_old[0]), .Y(\un18_next_int_m[0] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I249_Y (.A(I210_un1_Y), .B(
        ADD_26x26_fast_I210_Y_1), .C(ADD_26x26_fast_I249_Y_0), .Y(
        \un1_integ[19] ));
    GND GND_i (.Y(GND));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I146_un1_Y (.A(N470), .B(N477), 
        .Y(I146_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I104_un1_Y (.A(N426), .B(N423), 
        .Y(I104_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I6_P0N (.A(\un1_next_int[6] ), .B(
        integral[6]), .Y(N336));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I1_G0N (.A(\integ[1]_net_1 ), 
        .B(\un1_next_int[1] ), .Y(N320));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I107_Y (.A(N425), .B(N429), .Y(
        N478));
    NOR3B \state_RNI3F2A1[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[1] ), .Y(\un2_next_int_m[1] ));
    XNOR2 inf_abs1_a_1_I_9 (.A(sr_old[3]), .B(N_11), .Y(
        \inf_abs1_a_1[3] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I38_Y (.A(integral[17]), .B(
        integral[18]), .C(\un1_next_int_0_iv_0[13] ), .Y(N406));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I209_un1_Y_0 (.A(N543), .B(N512)
        , .Y(ADD_26x26_fast_I209_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_3 (.A(N504), .B(N519), .C(
        ADD_26x26_fast_I205_Y_2), .Y(ADD_26x26_fast_I205_Y_3));
    AX1D un1_integ_0_0_ADD_26x26_fast_I255_Y (.A(I204_un1_Y), .B(
        ADD_26x26_fast_I204_Y_3), .C(ADD_26x26_fast_I255_Y_0), .Y(
        \un1_integ[25] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I204_Y_0 (.A(integral[24]), .B(
        integral[23]), .C(\un1_next_int_0_iv[13] ), .Y(
        ADD_26x26_fast_I204_Y_0));
    MX2 \inf_abs0[4]  (.A(sr_new[4]), .B(\inf_abs0_a_0[4] ), .S(
        sr_new_0_0), .Y(\inf_abs0[4]_net_1 ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I243_Y (.A(N525), .B(I190_un1_Y), 
        .C(ADD_26x26_fast_I243_Y_0), .Y(\un1_integ[13] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I69_Y (.A(N324), .B(N327), .Y(
        N437));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I62_Y (.A(N332), .B(integral[6]), 
        .C(\un1_next_int[6] ), .Y(N430));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I193_un1_Y (.A(N478), .B(N486), 
        .C(N493), .Y(I193_un1_Y));
    NOR2B \state_RNIRPLN[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), .Y(
        next_int_0_sqmuxa_1));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I153_Y (.A(N484), .B(N476), .Y(
        N530));
    XNOR2 inf_abs0_a_0_I_7 (.A(sr_new[2]), .B(N_12), .Y(
        \inf_abs0_a_0[2] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I7_G0N (.A(\un2_next_int_m[7] ), 
        .B(\un1_next_int_iv_1[7] ), .C(integral[7]), .Y(N338));
    OA1A un1_integ_0_0_ADD_26x26_fast_I49_Y (.A(
        \un1_next_int_0_iv[13] ), .B(integral[13]), .C(N354), .Y(N417));
    OA1B un1_integ_0_0_ADD_26x26_fast_I42_Y (.A(integral[15]), .B(
        integral[16]), .C(\un1_next_int_0_iv_0[13] ), .Y(N410));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I145_Y (.A(N468), .B(N476), .Y(
        N522));
    MX2 \inf_abs1[4]  (.A(sr_old[4]), .B(\inf_abs1_a_1[4] ), .S(
        sr_old[12]), .Y(\inf_abs1[4]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I10_P0N (.A(integral[10]), .B(
        \un1_next_int[10] ), .Y(N348));
    OR2 un1_integ_0_0_ADD_26x26_fast_I1_P0N (.A(\integ[1]_net_1 ), .B(
        \un1_next_int[1] ), .Y(N321));
    OR3 \state_RNIM6V34[1]  (.A(\inf_abs1_m[3] ), .B(
        \un18_next_int_m[3] ), .C(\inf_abs0_m[3] ), .Y(
        \un1_next_int_iv_1[3] ));
    NOR3A inf_abs0_a_0_I_13 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .C(
        sr_new[4]), .Y(N_9_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I141_Y (.A(N419), .B(N423), .C(
        N464), .Y(N518));
    NOR2B \state_RNI42953_0[0]  (.A(\inf_abs0[11]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[11] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I93_Y (.A(N411), .B(N415), .Y(
        N464));
    AO1B un1_integ_0_0_ADD_26x26_fast_I37_Y (.A(integral[19]), .B(
        integral[18]), .C(\un1_next_int_0_iv_0[13] ), .Y(N405));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I0_G0N (.A(\integ[0]_net_1 ), 
        .B(N_3), .Y(N317));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I73_Y (.A(N318), .B(N321), .Y(
        N441));
    OA1 un1_integ_0_0_ADD_26x26_fast_I59_Y (.A(integral[8]), .B(
        \un1_next_int[8] ), .C(N339), .Y(N427));
    AO1 un1_integ_0_0_ADD_26x26_fast_I52_Y (.A(N347), .B(N351), .C(
        N350), .Y(N420));
    NOR2A \state_RNO[1]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 ), 
        .Y(\state_RNO_2[1] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I34_Y (.A(integral[20]), .B(
        integral[19]), .C(\un1_next_int_0_iv_0[13] ), .Y(N402));
    AX1D un1_integ_0_0_ADD_26x26_fast_I236_Y (.A(N485), .B(I161_un1_Y), 
        .C(ADD_26x26_fast_I236_Y_0), .Y(\un1_integ[6] ));
    NOR3C \state_RNIT4441[1]  (.A(sr_old[0]), .B(\state[1]_net_1 ), .C(
        sr_old[12]), .Y(\inf_abs1_m[0] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_1 (.A(N397), .B(N400), .C(
        ADD_26x26_fast_I205_Y_0), .Y(ADD_26x26_fast_I205_Y_1));
    OR2 un1_integ_0_0_ADD_26x26_fast_I150_Y (.A(I150_un1_Y), .B(N473), 
        .Y(N527));
    DFN1E0C0 \integ[0]  (.D(\un1_integ[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(\integ[0]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I120_Y (.A(I120_un1_Y), .B(N438), 
        .Y(N491));
    OR2 un1_integ_0_0_ADD_26x26_fast_I104_Y (.A(I104_un1_Y), .B(N422), 
        .Y(N475));
    VCC VCC_i (.Y(VCC));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I129_Y (.A(N452), .B(N460), .Y(
        N506));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I113_Y (.A(N431), .B(N435), .Y(
        N484));
    XNOR2 inf_abs0_a_0_I_28 (.A(sr_new[10]), .B(N_4_0), .Y(
        \inf_abs0_a_0[10] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I89_Y (.A(N407), .B(N411), .Y(
        N460));
    AO1 un1_integ_0_0_ADD_26x26_fast_I68_Y (.A(N323), .B(N327), .C(
        N326), .Y(N436));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_0 (.A(N462), .B(N469), .C(
        N461), .Y(ADD_26x26_fast_I211_Y_0));
    DFN1E0C0 \integ[4]  (.D(\un1_integ[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(\integ[4]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I108_Y (.A(N430), .B(N427), .C(
        N426), .Y(N479));
    NOR2B \state_RNIFOUS2[0]  (.A(\inf_abs0[6]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[6] ));
    NOR3 inf_abs1_a_1_I_18 (.A(sr_old[4]), .B(sr_old[3]), .C(sr_old[5])
        , .Y(\DWACT_FINC_E[2] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I3_G0N (.A(\integ[3]_net_1 ), 
        .B(\un1_next_int[3] ), .Y(N326));
    AO13 un1_integ_0_0_ADD_26x26_fast_I48_Y (.A(integral[13]), .B(N353)
        , .C(\un1_next_int_0_iv[13] ), .Y(N416));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I195_un1_Y (.A(N482), .B(N490), 
        .C(\state_RNICBRB4[0]_net_1 ), .Y(I195_un1_Y));
    DFN1E0C0 \integ[3]  (.D(\un1_integ[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(\integ[3]_net_1 ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I252_Y (.A(I174_un1_Y), .B(
        ADD_26x26_fast_I207_Y_2), .C(ADD_26x26_fast_I252_Y_0), .Y(
        \un1_integ[22] ));
    DFN1E0C0 \integ[6]  (.D(\un1_integ[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(integral[6]));
    XNOR2 inf_abs0_a_0_I_14 (.A(sr_new[5]), .B(N_9_0), .Y(
        \inf_abs0_a_0[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_1 (.A(N529), .B(N514), .C(
        ADD_26x26_fast_I210_Y_0), .Y(ADD_26x26_fast_I210_Y_1));
    AND3 inf_abs0_a_0_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[5] ), .Y(
        \DWACT_FINC_E[6] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y (.A(N533), .B(I194_un1_Y), 
        .C(ADD_26x26_fast_I239_Y_0), .Y(\un1_integ[9] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I106_un1_Y (.A(N428), .B(N425), 
        .Y(I106_un1_Y));
    NOR3A \state_RNI6E441[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .C(sr_old[9]), .Y(\un18_next_int_m[9] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_0 (.A(N402), .B(N399), .C(
        N398), .Y(ADD_26x26_fast_I206_Y_0));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I58_Y (.A(N338), .B(integral[8]), 
        .C(\un1_next_int[8] ), .Y(N426));
    OA1 un1_integ_0_0_ADD_26x26_fast_I67_Y (.A(\un1_next_int[4] ), .B(
        \integ[4]_net_1 ), .C(N327), .Y(N435));
    XNOR2 inf_abs0_a_0_I_12 (.A(sr_new[4]), .B(N_10), .Y(
        \inf_abs0_a_0[4] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I253_Y_0 (.A(integral[23]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I253_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I157_Y (.A(N488), .B(N480), .Y(
        N534));
    OR2 un1_integ_0_0_ADD_26x26_fast_I64_Y (.A(I64_un1_Y), .B(N332), 
        .Y(N432));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I204_un1_Y_0 (.A(N502), .B(N518)
        , .Y(ADD_26x26_fast_I204_un1_Y_0));
    NOR3B \state_RNIKQOR2[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[7] ), .Y(\un2_next_int_m[7] ));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I212_un1_Y (.A(N534), .B(N442), 
        .C(N518), .Y(I212_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I127_Y (.A(N458), .B(N450), .Y(
        N504));
    OR2 un1_integ_0_0_ADD_26x26_fast_I110_Y (.A(I110_un1_Y), .B(N428), 
        .Y(N481));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I211_un1_Y_0 (.A(N478), .B(N486)
        , .C(N493), .Y(ADD_26x26_fast_I211_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I90_Y (.A(N409), .B(N412), .C(
        N408), .Y(N461));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I233_Y (.A(
        ADD_26x26_fast_I233_Y_0), .B(N491), .Y(\un1_integ[3] ));
    NOR3A inf_abs0_a_0_I_31 (.A(\DWACT_FINC_E[6] ), .B(sr_new[9]), .C(
        sr_new[10]), .Y(N_3_1));
    AO1B un1_integ_0_0_ADD_26x26_fast_I47_Y (.A(integral[13]), .B(
        integral[14]), .C(\un1_next_int_0_iv[13] ), .Y(N415));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I119_Y (.A(N441), .B(N437), .Y(
        N490));
    AO1 un1_integ_0_0_ADD_26x26_fast_I70_Y (.A(N320), .B(N324), .C(
        N323), .Y(N438));
    NOR3A \state_RNI4C441[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .C(sr_old[7]), .Y(\un18_next_int_m[7] ));
    DFN1E0C0 \integ[5]  (.D(\un1_integ[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(\integ[5]_net_1 ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I44_Y (.A(integral[14]), .B(
        integral[15]), .C(\un1_next_int_0_iv_0[13] ), .Y(N412));
    AX1D un1_integ_0_0_ADD_26x26_fast_I245_Y (.A(N521), .B(I188_un1_Y), 
        .C(ADD_26x26_fast_I245_Y_0), .Y(\un1_integ[15] ));
    NOR2 \state_RNIB7PP_0[0]  (.A(\state[1]_net_1 ), .B(
        \state[0]_net_1 ), .Y(N_46_1_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I95_Y (.A(N413), .B(N417), .Y(
        N466));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y_0 (.A(\un2_next_int_m[9] )
        , .B(\un1_next_int_iv_1[9] ), .C(integral[9]), .Y(
        ADD_26x26_fast_I239_Y_0));
    DFN1E0C0 \integ[2]  (.D(\un1_integ[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(\integ[2]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I135_Y (.A(N458), .B(N466), .Y(
        N512));
    OR2 un1_integ_0_0_ADD_26x26_fast_I88_Y (.A(N410), .B(N406), .Y(
        N459));
    AX1D un1_integ_0_0_ADD_26x26_fast_I247_Y (.A(I212_un1_Y), .B(
        ADD_26x26_fast_I212_Y_0), .C(ADD_26x26_fast_I247_Y_0), .Y(
        \un1_integ[17] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I237_Y_0 (.A(\un2_next_int_m[7] )
        , .B(\un1_next_int_iv_1[7] ), .C(integral[7]), .Y(
        ADD_26x26_fast_I237_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I143_Y (.A(N466), .B(N474), .Y(
        N520));
    OR3 \state_RNIJQ1A3[0]  (.A(\inf_abs1_m[0] ), .B(
        \un18_next_int_m[0] ), .C(\inf_abs0_m[0] ), .Y(
        \un1_next_int_iv_1[0] ));
    NOR2B \state_RNIDIBM[0]  (.A(sr_new[3]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[3] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I57_Y (.A(integral[8]), .B(
        \un1_next_int[8] ), .C(N345), .Y(N425));
    OA1 un1_integ_0_0_ADD_26x26_fast_I186_un1_Y (.A(N481), .B(
        I158_un1_Y), .C(N520), .Y(I186_un1_Y));
    NOR3 inf_abs0_a_0_I_29 (.A(sr_new[7]), .B(sr_new[6]), .C(sr_new[8])
        , .Y(\DWACT_FINC_E_0[5] ));
    OR3 \state_RNISHPL5[1]  (.A(\inf_abs0_m[7] ), .B(
        \un18_next_int_m[7] ), .C(\inf_abs1_m[7] ), .Y(
        \un1_next_int_iv_1[7] ));
    DFN1E0C0 \integ[23]  (.D(\un1_integ[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[23]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_2 (.A(
        ADD_26x26_fast_I206_un1_Y_0), .B(N522), .C(
        ADD_26x26_fast_I206_Y_1), .Y(ADD_26x26_fast_I206_Y_2));
    AO1 un1_integ_0_0_ADD_26x26_fast_I54_Y (.A(N344), .B(N348), .C(
        N347), .Y(N422));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I131_Y (.A(N454), .B(N462), .Y(
        N508));
    XNOR2 inf_abs0_a_0_I_26 (.A(sr_new[9]), .B(N_5), .Y(
        \inf_abs0_a_0[9] ));
    NOR3B inf_abs1_a_1_I_19 (.A(\DWACT_FINC_E[2] ), .B(
        \DWACT_FINC_E_0[0] ), .C(sr_old[6]), .Y(N_7));
    OR2 \state_RNISBO51[1]  (.A(next_int_1_sqmuxa), .B(
        next_int_0_sqmuxa_1), .Y(\un1_next_int_0_iv_0[13] ));
    NOR3B inf_abs1_a_1_I_16 (.A(\DWACT_FINC_E[1] ), .B(
        \DWACT_FINC_E_0[0] ), .C(sr_old[5]), .Y(N_8));
    NOR3B \state_RNI16VO3[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[8]_net_1 ), .Y(\un2_next_int_m[8] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I254_Y (.A(I205_un1_Y), .B(
        ADD_26x26_fast_I205_Y_3), .C(ADD_26x26_fast_I254_Y_0), .Y(
        \un1_integ[24] ));
    DFN1E0C0 \integ[19]  (.D(\un1_integ[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[19]));
    NOR2 inf_abs0_a_0_I_15 (.A(sr_new[3]), .B(sr_new[4]), .Y(
        \DWACT_FINC_E_0[1] ));
    MX2 \inf_abs1[8]  (.A(sr_old[8]), .B(\inf_abs1_a_1[8] ), .S(
        sr_old[12]), .Y(\inf_abs1[8]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I161_un1_Y (.A(N486), .B(N493), 
        .Y(I161_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I117_Y (.A(N439), .B(N435), .Y(
        N488));
    DFN1E0C0 \integ[17]  (.D(\un1_integ[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[17]));
    XOR2 inf_abs0_a_0_I_5 (.A(sr_new[0]), .B(sr_new[1]), .Y(
        \inf_abs0_a_0[1] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I33_Y (.A(integral[20]), .B(
        integral[21]), .C(\un1_next_int_0_iv_0[13] ), .Y(N401));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I255_Y_0 (.A(integral[25]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I255_Y_0));
    DFN1E0C0 \integ[14]  (.D(\un1_integ[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[14]));
    XNOR2 inf_abs0_a_0_I_17 (.A(sr_new[6]), .B(N_8_0), .Y(
        \inf_abs0_a_0[6] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I87_Y (.A(N405), .B(N409), .Y(
        N458));
    AO1B un1_integ_0_0_ADD_26x26_fast_I29_Y (.A(integral[23]), .B(
        integral[22]), .C(\un1_next_int_0_iv_0[13] ), .Y(N397));
    OR2 un1_integ_0_0_ADD_26x26_fast_I84_Y (.A(N406), .B(N402), .Y(
        N455));
    AO1 un1_integ_0_0_ADD_26x26_fast_I154_Y (.A(N485), .B(N478), .C(
        N477), .Y(N531));
    MX2 \inf_abs1[11]  (.A(sr_old[11]), .B(\inf_abs1_a_1[11] ), .S(
        sr_old[12]), .Y(\inf_abs1[11]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I11_G0N (.A(integral[11]), .B(
        \state_RNIKDT9C[0]_net_1 ), .Y(N350));
    OR2 \state_RNIGLJU5[0]  (.A(\un1_next_int_iv_1[3] ), .B(
        \un2_next_int_m[3] ), .Y(\un1_next_int[3] ));
    XA1A \state_RNIRJ264[1]  (.A(sr_old[12]), .B(\inf_abs1[6]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[6] ));
    MX2 \inf_abs1[2]  (.A(sr_old[2]), .B(\inf_abs1_a_1[2] ), .S(
        sr_old[12]), .Y(\inf_abs1[2]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I140_Y (.A(N471), .B(N464), .C(
        N463), .Y(N517));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I149_Y (.A(N419), .B(N423), .C(
        N480), .Y(N526));
    OR3 \state_RNI86EBA[0]  (.A(\inf_abs0_m[6] ), .B(
        \un1_next_int_iv_0[6] ), .C(\un2_next_int_m[6] ), .Y(
        \un1_next_int[6] ));
    NOR3B \state_RNIPGP11_0[0]  (.A(\state[0]_net_1 ), .B(sr_new_0_0), 
        .C(sr_new[0]), .Y(\un2_next_int_m[0] ));
    NOR2B \state_RNII4HD3[0]  (.A(\inf_abs0[8]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[8] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I249_Y_0 (.A(integral[19]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I249_Y_0));
    INV \integ_RNIH9BD[24]  (.A(integral[24]), .Y(integral_i[24]));
    DFN1E0C0 \integ[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[25]));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I247_Y_0 (.A(integral[17]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I247_Y_0));
    NOR3B \state_RNI4E872[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[2]_net_1 ), .Y(\un2_next_int_m[2] ));
    MX2 \inf_abs1[6]  (.A(sr_old[6]), .B(\inf_abs1_a_1[6] ), .S(
        sr_old[12]), .Y(\inf_abs1[6]_net_1 ));
    NOR3 inf_abs0_a_0_I_33 (.A(sr_new[10]), .B(sr_new[9]), .C(
        sr_new[11]), .Y(\DWACT_FINC_E[7] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y_0 (.A(\integ[0]_net_1 ), 
        .B(N_3), .Y(ADD_26x26_fast_I230_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I64_un1_Y (.A(N329), .B(N333), 
        .Y(I64_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I242_Y (.A(N527), .B(I191_un1_Y), 
        .C(ADD_26x26_fast_I242_Y_0), .Y(\un1_integ[12] ));
    XNOR2 inf_abs0_a_0_I_20 (.A(sr_new[7]), .B(N_7_0), .Y(
        \inf_abs0_a_0[7] ));
    DFN1E0C0 \integ[11]  (.D(\un1_integ[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[11]));
    MX2 \inf_abs0[8]  (.A(sr_new[8]), .B(\inf_abs0_a_0[8] ), .S(
        sr_new_0_0), .Y(\inf_abs0[8]_net_1 ));
    DFN1E0C0 \integ[16]  (.D(\un1_integ[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[16]));
    XNOR2 inf_abs1_a_1_I_28 (.A(sr_old[10]), .B(N_4), .Y(
        \inf_abs1_a_1[10] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I211_Y_1 (.A(
        ADD_26x26_fast_I211_un1_Y_0), .B(N531), .C(
        ADD_26x26_fast_I211_Y_1_0), .Y(ADD_26x26_fast_I211_Y_1));
    NOR3 inf_abs1_a_1_I_10 (.A(sr_old[1]), .B(sr_old[0]), .C(sr_old[2])
        , .Y(\DWACT_FINC_E_0[0] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I254_Y_0 (.A(integral[24]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I254_Y_0));
    OR3 un1_integ_0_0_ADD_26x26_fast_I163_Y (.A(N436), .B(I118_un1_Y), 
        .C(I163_un1_Y), .Y(N543));
    MX2B un1_next_int_0_sqmuxa_0__m2 (.A(sr_new_1_0), .B(sr_old[12]), 
        .S(\state[1]_net_1 ), .Y(N_3));
    AO1 un1_integ_0_0_ADD_26x26_fast_I96_Y (.A(N418), .B(N415), .C(
        N414), .Y(N467));
    MX2 \inf_abs0[10]  (.A(sr_new[10]), .B(\inf_abs0_a_0[10] ), .S(
        sr_new_1_0), .Y(\inf_abs0[10]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I2_G0N (.A(\integ[2]_net_1 ), 
        .B(\un1_next_int[2] ), .Y(N323));
    AO1 un1_integ_0_0_ADD_26x26_fast_I114_Y (.A(N436), .B(N433), .C(
        N432), .Y(N485));
    OA1 un1_integ_0_0_ADD_26x26_fast_I189_un1_Y (.A(N485), .B(
        I161_un1_Y), .C(N524), .Y(I189_un1_Y));
    MX2 \inf_abs1[1]  (.A(sr_old[1]), .B(\inf_abs1_a_1[1] ), .S(
        sr_old[12]), .Y(\inf_abs1[1]_net_1 ));
    NOR2 inf_abs0_a_0_I_21 (.A(sr_new[6]), .B(sr_new[7]), .Y(
        \DWACT_FINC_E_0[3] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I147_Y (.A(N470), .B(N478), .Y(
        N524));
    DFN1E0C0 \integ[9]  (.D(\un1_integ[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(integral[9]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I242_Y_0 (.A(
        \un2_next_int_m[12] ), .B(\un1_next_int_iv_0[12] ), .C(
        integral[12]), .Y(ADD_26x26_fast_I242_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I235_Y (.A(N487), .B(I162_un1_Y), 
        .C(ADD_26x26_fast_I235_Y_0), .Y(\un1_integ[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I212_Y_0 (.A(N533), .B(N518), .C(
        N517), .Y(ADD_26x26_fast_I212_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I63_Y (.A(N333), .B(N336), .Y(
        N431));
    NOR2A inf_abs1_a_1_I_11 (.A(\DWACT_FINC_E_0[0] ), .B(sr_old[3]), 
        .Y(N_10_0));
    OR3 \state_RNIPICH8[0]  (.A(\inf_abs0_m[4] ), .B(
        \un1_next_int_iv_0[4] ), .C(\un2_next_int_m[4] ), .Y(
        \un1_next_int[4] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I237_Y (.A(N483), .B(I160_un1_Y), 
        .C(ADD_26x26_fast_I237_Y_0), .Y(\un1_integ[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I133_Y (.A(N456), .B(N464), .Y(
        N510));
    NOR3B \state_RNI42953[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[11]_net_1 ), .Y(\un2_next_int_m[11] ));
    NOR2B \state_RNIGGCC2[0]  (.A(\inf_abs0[4]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[4] ));
    MX2 \inf_abs0[2]  (.A(sr_new[2]), .B(\inf_abs0_a_0[2] ), .S(
        sr_new_0_0), .Y(\inf_abs0[2]_net_1 ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I30_Y (.A(integral[22]), .B(
        integral[21]), .C(\un1_next_int_0_iv_0[13] ), .Y(N398));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I160_un1_Y (.A(N484), .B(N491), 
        .Y(I160_un1_Y));
    DFN1E0C0 \integ[22]  (.D(\un1_integ[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[22]));
    NOR3 inf_abs1_a_1_I_8 (.A(sr_old[1]), .B(sr_old[0]), .C(sr_old[2]), 
        .Y(N_11));
    AO1B un1_integ_0_0_ADD_26x26_fast_I43_Y (.A(integral[15]), .B(
        integral[16]), .C(\un1_next_int_0_iv_0[13] ), .Y(N411));
    NOR3B \state_RNIVHQN2[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[4]_net_1 ), .Y(\un2_next_int_m[4] ));
    OR3 \state_RNI7ASS4[1]  (.A(\inf_abs0_m[5] ), .B(
        \un18_next_int_m[5] ), .C(\inf_abs1_m[5] ), .Y(
        \un1_next_int_iv_1[5] ));
    DFN1E0C0 \integ_0[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral_0_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I192_Y (.A(N530), .B(N491), .C(
        N529), .Y(N649));
    DFN1E0C0 \integ[1]  (.D(\un1_integ[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(\integ[1]_net_1 ));
    OR3 \state_RNIKDT9C[0]  (.A(\inf_abs0_m[11] ), .B(
        \un1_next_int_iv_0[11] ), .C(\un2_next_int_m[11] ), .Y(
        \state_RNIKDT9C[0]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I35_Y (.A(integral[19]), .B(
        integral[20]), .C(\un1_next_int_0_iv_0[13] ), .Y(N403));
    NOR2B inf_abs0_a_0_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_2));
    INV \integ_RNIIABD[25]  (.A(integral[25]), .Y(integral_i[25]));
    OR2 un1_integ_0_0_ADD_26x26_fast_I204_Y_1 (.A(
        ADD_26x26_fast_I204_Y_0), .B(N398), .Y(ADD_26x26_fast_I204_Y_1)
        );
    NOR2B un1_integ_0_0_ADD_26x26_fast_I53_Y (.A(N351), .B(N348), .Y(
        N421));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I91_Y (.A(N409), .B(N413), .Y(
        N462));
    AX1D un1_integ_0_0_ADD_26x26_fast_I250_Y (.A(I178_un1_Y), .B(
        ADD_26x26_fast_I209_Y_1), .C(ADD_26x26_fast_I250_Y_0), .Y(
        \un1_integ[20] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I240_Y_0 (.A(integral[10]), .B(
        \un1_next_int[10] ), .Y(ADD_26x26_fast_I240_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I60_un1_Y (.A(integral[6]), .B(
        \un1_next_int[6] ), .C(N339), .Y(I60_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_0 (.A(N467), .B(N460), .C(
        N459), .Y(ADD_26x26_fast_I210_Y_0));
    NOR2B \state_RNIFKBM[0]  (.A(sr_new[5]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[5] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I71_Y (.A(N321), .B(N324), .Y(
        N439));
    DFN1E0C0 \integ[20]  (.D(\un1_integ[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[20]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I244_Y (.A(N523), .B(I189_un1_Y), 
        .C(ADD_26x26_fast_I244_Y_0), .Y(\un1_integ[14] ));
    NOR2A \state_RNI1I2E[0]  (.A(\state[0]_net_1 ), .B(sr_new[12]), .Y(
        next_int_1_sqmuxa));
    NOR3 inf_abs1_a_1_I_29 (.A(sr_old[8]), .B(sr_old[7]), .C(sr_old[6])
        , .Y(\DWACT_FINC_E[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_1 (.A(N454), .B(N461), .C(
        ADD_26x26_fast_I207_Y_0), .Y(ADD_26x26_fast_I207_Y_1));
    OR2 un1_integ_0_0_ADD_26x26_fast_I106_Y (.A(I106_un1_Y), .B(N424), 
        .Y(N477));
    XNOR2 inf_abs0_a_0_I_32 (.A(sr_new[11]), .B(N_3_1), .Y(
        \inf_abs0_a_0[11] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_1 (.A(
        ADD_26x26_fast_I208_un1_Y_0), .B(N526), .C(
        ADD_26x26_fast_I208_Y_0), .Y(ADD_26x26_fast_I208_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I102_Y (.A(N424), .B(N421), .C(
        N420), .Y(N473));
    NOR2B \state_RNIMBC23[1]  (.A(\inf_abs1_a_1[5] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[5] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I251_Y (.A(I176_un1_Y), .B(
        ADD_26x26_fast_I208_Y_1), .C(ADD_26x26_fast_I251_Y_0), .Y(
        \un1_integ[21] ));
    XNOR2 inf_abs1_a_1_I_26 (.A(sr_old[9]), .B(N_5_0), .Y(
        \inf_abs1_a_1[9] ));
    DFN1E0C0 \integ[18]  (.D(\un1_integ[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[18]));
    OR2 un1_integ_0_0_ADD_26x26_fast_I144_Y (.A(I144_un1_Y), .B(N467), 
        .Y(N521));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I83_Y (.A(N405), .B(N401), .Y(
        N454));
    NOR2B \state_RNI83343_0[0]  (.A(\inf_abs0[10]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[10] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_0 (.A(N458), .B(N465), .C(
        N457), .Y(ADD_26x26_fast_I209_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_0 (.A(N401), .B(N404), .C(
        N400), .Y(ADD_26x26_fast_I207_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I148_Y (.A(I148_un1_Y), .B(N471), 
        .Y(N525));
    XA1A \state_RNIO2Q72[1]  (.A(sr_old[12]), .B(\inf_abs1[1]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[1] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I60_Y (.A(I60_un1_Y), .B(N338), 
        .Y(N428));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I232_Y (.A(\un1_next_int[2] ), 
        .B(\integ[2]_net_1 ), .C(N493), .Y(\un1_integ[2] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I204_Y_2 (.A(N455), .B(N448), .C(
        ADD_26x26_fast_I204_Y_1), .Y(ADD_26x26_fast_I204_Y_2));
    DFN1C0 \state[1]  (.D(\state_RNO_2[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[1]_net_1 ));
    XNOR2 inf_abs0_a_0_I_23 (.A(sr_new[8]), .B(N_6_0), .Y(
        \inf_abs0_a_0[8] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I118_un1_Y (.A(N440), .B(N437), 
        .Y(I118_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I110_un1_Y (.A(N432), .B(N429), 
        .Y(I110_un1_Y));
    NOR3A inf_abs1_a_1_I_13 (.A(\DWACT_FINC_E_0[0] ), .B(sr_old[3]), 
        .C(sr_old[4]), .Y(N_9));
    OA1 un1_integ_0_0_ADD_26x26_fast_I9_G0N (.A(\un2_next_int_m[9] ), 
        .B(\un1_next_int_iv_1[9] ), .C(integral[9]), .Y(N344));
    OA1B un1_integ_0_0_ADD_26x26_fast_I40_Y (.A(integral[17]), .B(
        integral[16]), .C(\un1_next_int_0_iv_0[13] ), .Y(N408));
    OA1 un1_integ_0_0_ADD_26x26_fast_I65_Y (.A(\un1_next_int[4] ), .B(
        \integ[4]_net_1 ), .C(N333), .Y(N433));
    XA1A \state_RNIGRVU4[1]  (.A(sr_old[12]), .B(\inf_abs1[8]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[8] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I207_un1_Y_0 (.A(N485), .B(
        I161_un1_Y), .C(N508), .Y(ADD_26x26_fast_I207_un1_Y_0));
    NOR3B \state_RNIPUE43[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[12] ), .Y(\un2_next_int_m[12] ));
    NOR3 inf_abs0_a_0_I_8 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2]), 
        .Y(N_11_0));
    AND3 inf_abs1_a_1_I_30 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E_0[6] ));
    XNOR2 inf_abs0_a_0_I_35 (.A(sr_new[12]), .B(N_2), .Y(
        \inf_abs0_a_0[12] ));
    NOR2B \state_RNI7F9R3[1]  (.A(\inf_abs1_a_1[7] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I178_un1_Y (.A(N512), .B(N527), 
        .Y(I178_un1_Y));
    AO1B un1_integ_0_0_ADD_26x26_fast_I45_Y (.A(integral[15]), .B(
        integral[14]), .C(\un1_next_int_0_iv_0[13] ), .Y(N413));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I137_Y (.A(N468), .B(N460), .Y(
        N514));
    NOR3B \state_RNIQEKQ1[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[3] ), .Y(\un2_next_int_m[3] ));
    XNOR2 inf_abs0_a_0_I_9 (.A(sr_new[3]), .B(N_11_0), .Y(
        \inf_abs0_a_0[3] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I3_P0N (.A(\integ[3]_net_1 ), .B(
        \un1_next_int[3] ), .Y(N327));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I233_Y_0 (.A(\integ[3]_net_1 ), 
        .B(\un1_next_int[3] ), .Y(ADD_26x26_fast_I233_Y_0));
    NOR2B \state_RNO[0]  (.A(N_46_1), .B(calc_int), .Y(
        \state_RNO_1[0] ));
    NOR3A \state_RNI2A441[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .C(sr_old[5]), .Y(\un18_next_int_m[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I50_Y (.A(N350), .B(N354), .C(
        N353), .Y(N418));
    AO1 un1_integ_0_0_ADD_26x26_fast_I204_Y_3 (.A(N517), .B(N502), .C(
        ADD_26x26_fast_I204_Y_2), .Y(ADD_26x26_fast_I204_Y_3));
    XNOR2 inf_abs1_a_1_I_20 (.A(sr_old[7]), .B(N_7), .Y(
        \inf_abs1_a_1[7] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I36_Y (.A(integral[18]), .B(
        integral[19]), .C(\un1_next_int_0_iv_0[13] ), .Y(N404));
    NOR3A inf_abs1_a_1_I_31 (.A(\DWACT_FINC_E_0[6] ), .B(sr_old[9]), 
        .C(sr_old[10]), .Y(N_3_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I0_P0N (.A(\integ[0]_net_1 ), .B(
        N_3), .Y(N318));
    NOR2 inf_abs1_a_1_I_6 (.A(sr_old[0]), .B(sr_old[1]), .Y(N_12_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I77_Y_0 (.A(integral[23]), .B(
        integral[24]), .C(\un1_next_int_0_iv[13] ), .Y(
        ADD_26x26_fast_I77_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I55_Y (.A(N345), .B(N348), .Y(
        N423));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I205_un1_Y (.A(N520), .B(N504), 
        .C(N658), .Y(I205_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I163_un1_Y (.A(N490), .B(
        \state_RNICBRB4[0]_net_1 ), .Y(I163_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I120_un1_Y (.A(N439), .B(N442), 
        .Y(I120_un1_Y));
    OR3 \state_RNI36G5C[0]  (.A(\inf_abs0_m[8] ), .B(
        \un1_next_int_iv_0[8] ), .C(\un2_next_int_m[8] ), .Y(
        \un1_next_int[8] ));
    NOR2 inf_abs1_a_1_I_21 (.A(sr_old[7]), .B(sr_old[6]), .Y(
        \DWACT_FINC_E[3] ));
    NOR2B \state_RNIJOBM[0]  (.A(sr_new[9]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[9] ));
    NOR2B \state_RNI9CF92[1]  (.A(\inf_abs1_a_1[3] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[3] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_1 (.A(N459), .B(N452), .C(
        ADD_26x26_fast_I206_Y_0), .Y(ADD_26x26_fast_I206_Y_1));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I5_G0N (.A(\integ[5]_net_1 ), 
        .B(\un1_next_int[5] ), .Y(N332));
    AND3 inf_abs0_a_0_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(
        \DWACT_FINC_E[4] ));
    OR3 \state_RNIMBBN6[0]  (.A(\inf_abs0_m[2] ), .B(
        \un1_next_int_iv_0[2] ), .C(\un2_next_int_m[2] ), .Y(
        \un1_next_int[2] ));
    DFN1E0C0 \integ[7]  (.D(\un1_integ[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(integral[7]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_2 (.A(
        ADD_26x26_fast_I207_un1_Y_0), .B(N524), .C(
        ADD_26x26_fast_I207_Y_1), .Y(ADD_26x26_fast_I207_Y_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I4_G0N (.A(\integ[4]_net_1 ), 
        .B(\un1_next_int[4] ), .Y(N329));
    OR3 un1_integ_0_0_ADD_26x26_fast_I195_Y (.A(N481), .B(I158_un1_Y), 
        .C(I195_un1_Y), .Y(N658));
    OA1 un1_integ_0_0_ADD_26x26_fast_I206_un1_Y_0 (.A(N483), .B(
        I160_un1_Y), .C(N506), .Y(ADD_26x26_fast_I206_un1_Y_0));
    XNOR2 inf_abs1_a_1_I_14 (.A(sr_old[5]), .B(N_9), .Y(
        \inf_abs1_a_1[5] ));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I234_Y (.A(\un1_next_int[4] ), 
        .B(\integ[4]_net_1 ), .C(N543), .Y(\un1_integ[4] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_2 (.A(N450), .B(N457), .C(
        ADD_26x26_fast_I205_Y_1), .Y(ADD_26x26_fast_I205_Y_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I174_un1_Y (.A(N508), .B(N523), 
        .Y(I174_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I162_un1_Y (.A(N488), .B(N442), 
        .Y(I162_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I240_Y (.A(N531), .B(I193_un1_Y), 
        .C(ADD_26x26_fast_I240_Y_0), .Y(\un1_integ[10] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I156_Y (.A(N487), .B(N480), .C(
        N479), .Y(N533));
    DFN1E0C0 \integ[8]  (.D(\un1_integ[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(integral[8]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I85_Y (.A(N407), .B(N403), .Y(
        N456));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I251_Y_0 (.A(integral[21]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I251_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I152_Y (.A(N483), .B(N476), .C(
        N475), .Y(N529));
    AND3 inf_abs0_a_0_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(N_6_0));
    OR3 un1_integ_0_0_ADD_26x26_fast_I9_P0N (.A(\un2_next_int_m[9] ), 
        .B(\un1_next_int_iv_1[9] ), .C(integral[9]), .Y(N345));
    OA1 un1_integ_0_0_ADD_26x26_fast_I208_un1_Y_0 (.A(N487), .B(
        I162_un1_Y), .C(N510), .Y(ADD_26x26_fast_I208_un1_Y_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I31_Y (.A(integral[21]), .B(
        integral[22]), .C(\un1_next_int_0_iv_0[13] ), .Y(N399));
    XNOR2 inf_abs1_a_1_I_12 (.A(sr_old[4]), .B(N_10_0), .Y(
        \inf_abs1_a_1[4] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I235_Y_0 (.A(\integ[5]_net_1 ), 
        .B(\un1_next_int[5] ), .Y(ADD_26x26_fast_I235_Y_0));
    NOR3B \state_RNIUPC83[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[6]_net_1 ), .Y(\un2_next_int_m[6] ));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I241_Y (.A(
        \state_RNIKDT9C[0]_net_1 ), .B(integral[11]), .C(N649), .Y(
        \un1_integ[11] ));
    NOR3 inf_abs0_a_0_I_18 (.A(sr_new[3]), .B(sr_new[5]), .C(sr_new[4])
        , .Y(\DWACT_FINC_E_0[2] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I11_P0N (.A(integral[11]), .B(
        \state_RNIKDT9C[0]_net_1 ), .Y(N351));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I243_Y_0 (.A(integral[13]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I243_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I105_Y (.A(N427), .B(N423), .Y(
        N476));
    OR2 \state_RNICBRB4[0]  (.A(\un1_next_int_iv_1[0] ), .B(
        \un2_next_int_m[0] ), .Y(\state_RNICBRB4[0]_net_1 ));
    OR3 \state_RNILTME6[1]  (.A(\inf_abs0_m[9] ), .B(
        \un18_next_int_m[9] ), .C(\inf_abs1_m[9] ), .Y(
        \un1_next_int_iv_1[9] ));
    MX2 \inf_abs0[11]  (.A(sr_new[11]), .B(\inf_abs0_a_0[11] ), .S(
        sr_new_1_0), .Y(\inf_abs0[11]_net_1 ));
    NOR3B \state_RNIPGP11[0]  (.A(\state[0]_net_1 ), .B(sr_new[0]), .C(
        sr_new_0_0), .Y(\inf_abs0_m[0] ));
    XA1A \state_RNIC9BV5[1]  (.A(sr_old[12]), .B(\inf_abs1[11]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[11] ));
    XOR2 inf_abs1_a_1_I_5 (.A(sr_old[0]), .B(sr_old[1]), .Y(
        \inf_abs1_a_1[1] ));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I66_Y (.A(N326), .B(
        \un1_next_int[4] ), .C(\integ[4]_net_1 ), .Y(N434));
    AX1D un1_integ_0_0_ADD_26x26_fast_I248_Y (.A(
        ADD_26x26_fast_I211_Y_1), .B(ADD_26x26_fast_I211_Y_0), .C(
        ADD_26x26_fast_I248_Y_0), .Y(\un1_integ[18] ));
    OR2 \state_RNI62884[0]  (.A(\un1_next_int_iv_1[1] ), .B(
        \un2_next_int_m[1] ), .Y(\un1_next_int[1] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I99_Y (.A(N417), .B(N421), .Y(
        N470));
    OR2 un1_integ_0_0_ADD_26x26_fast_I92_Y (.A(N414), .B(N410), .Y(
        N463));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I191_un1_Y (.A(N528), .B(N543), 
        .Y(I191_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I79_Y (.A(N397), .B(N401), .Y(
        N450));
    AO1 un1_integ_0_0_ADD_26x26_fast_I72_Y (.A(N317), .B(N321), .C(
        N320), .Y(N440));
    NOR3B \state_RNI83343[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[10]_net_1 ), .Y(\un2_next_int_m[10] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I46_Y (.A(integral[13]), .B(
        integral[14]), .C(\un1_next_int_0_iv_0[13] ), .Y(N414));
    NOR3 inf_abs1_a_1_I_33 (.A(sr_old[10]), .B(sr_old[9]), .C(
        sr_old[11]), .Y(\DWACT_FINC_E_0[7] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I116_Y (.A(N438), .B(N435), .C(
        N434), .Y(N487));
    AO1 un1_integ_0_0_ADD_26x26_fast_I112_Y (.A(N434), .B(N431), .C(
        N430), .Y(N483));
    NOR2A inf_abs0_a_0_I_25 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .Y(
        N_5));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I8_G0N (.A(\un1_next_int[8] ), 
        .B(integral[8]), .Y(N341));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I213_un1_Y_0 (.A(N482), .B(N490)
        , .C(\state_RNICBRB4[0]_net_1 ), .Y(
        ADD_26x26_fast_I213_un1_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I210_un1_Y (.A(N514), .B(N491), 
        .C(N530), .Y(I210_un1_Y));
    NOR3A inf_abs0_a_0_I_27 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .C(
        sr_new[9]), .Y(N_4_0));
    
endmodule


module error_calc_13s_12s_4_0(
       cur_error,
       LED_33_i_0,
       LED_33,
       average,
       calc_error,
       n_rst_c,
       clk_c
    );
output [12:0] cur_error;
input  LED_33_i_0;
input  [7:0] LED_33;
input  [6:2] average;
input  calc_error;
input  n_rst_c;
input  clk_c;

    wire N_40, N_38, GND, VCC;
    
    AX1B un2_diffreg_1_m37 (.A(LED_33[5]), .B(LED_33[6]), .C(LED_33[7])
        , .Y(N_38));
    DFN1E1C0 \diffreg[3]  (.D(average[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[3]));
    XNOR2 un2_diffreg_1_m39 (.A(LED_33[6]), .B(LED_33[5]), .Y(N_40));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \diffreg[7]  (.D(LED_33[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[7]));
    DFN1E1C0 \diffreg[1]  (.D(average[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[1]));
    DFN1E1C0 \diffreg[12]  (.D(N_38), .CLK(clk_c), .CLR(n_rst_c), .E(
        calc_error), .Q(cur_error[12]));
    DFN1E1C0 \diffreg[11]  (.D(N_40), .CLK(clk_c), .CLR(n_rst_c), .E(
        calc_error), .Q(cur_error[11]));
    GND GND_i (.Y(GND));
    DFN1E1C0 \diffreg[9]  (.D(LED_33[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[9]));
    DFN1E1C0 \diffreg[8]  (.D(LED_33[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[8]));
    DFN1E1C0 \diffreg[6]  (.D(LED_33[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[6]));
    DFN1E1C0 \diffreg[10]  (.D(LED_33_i_0), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[10]));
    DFN1E1C0 \diffreg[5]  (.D(LED_33[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[5]));
    DFN1E1C0 \diffreg[4]  (.D(average[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[4]));
    DFN1E1C0 \diffreg[2]  (.D(average[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[2]));
    DFN1E1C0 \diffreg[0]  (.D(average[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[0]));
    
endmodule


module derivative_calc_13s_4_0(
       derivative_0,
       sr_prev,
       sr_new,
       sr_new_1_0,
       deriv_enable,
       n_rst_c,
       clk_c
    );
output derivative_0;
input  [12:0] sr_prev;
input  [11:0] sr_new;
input  sr_new_1_0;
input  deriv_enable;
input  n_rst_c;
input  clk_c;

    wire SUB_13x13_medium_area_I49_Y_1, N208, N176, 
        SUB_13x13_medium_area_I49_Y_0, 
        SUB_13x13_medium_area_I26_un1_Y_0, 
        SUB_13x13_medium_area_I49_un1_Y_1, 
        SUB_13x13_medium_area_I49_un1_Y_0, N_15, 
        SUB_13x13_medium_area_I42_Y_1, N218, N180, 
        SUB_13x13_medium_area_I42_Y_0, 
        SUB_13x13_medium_area_I30_un1_Y_0, 
        SUB_13x13_medium_area_I42_un1_Y_1, N_9, N_7, 
        SUB_13x13_medium_area_I41_Y_0, 
        SUB_13x13_medium_area_I34_un1_Y_0, 
        SUB_13x13_medium_area_I41_un1_Y_0, N_5, 
        SUB_13x13_medium_area_I32_un1_Y_0, 
        SUB_13x13_medium_area_I28_un1_Y_0, N_24, N226, N204, N212, 
        N222, N185, N_21, N_13, GND, VCC;
    
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I34_un1_Y_0 (.A(
        sr_new[1]), .B(sr_prev[1]), .Y(
        SUB_13x13_medium_area_I34_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y_0 (.A(
        SUB_13x13_medium_area_I30_un1_Y_0), .B(sr_new[6]), .C(
        sr_prev[6]), .Y(SUB_13x13_medium_area_I42_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I15_S (.A(sr_prev[2]), 
        .B(sr_new[2]), .Y(N_5));
    OR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I36_Y (.A(sr_prev[0]), 
        .B(sr_new[0]), .Y(N185));
    XNOR3 un2_deriv_out_0_0_SUB_13x13_medium_area_I82_Y (.A(sr_new_1_0)
        , .B(sr_prev[12]), .C(N226), .Y(N_24));
    VCC VCC_i (.Y(VCC));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I64_Y (.A(N204), .B(
        sr_new[11]), .C(sr_prev[11]), .Y(N226));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I41_Y_0 (.A(
        SUB_13x13_medium_area_I34_un1_Y_0), .B(sr_new[2]), .C(
        sr_prev[2]), .Y(SUB_13x13_medium_area_I41_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I19_S (.A(sr_prev[6]), 
        .B(sr_new[6]), .Y(N_13));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I28_Y (.A(
        SUB_13x13_medium_area_I28_un1_Y_0), .B(sr_new[8]), .C(
        sr_prev[8]), .Y(N208));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y_1 (.A(N218), .B(
        N180), .C(SUB_13x13_medium_area_I42_Y_0), .Y(
        SUB_13x13_medium_area_I42_Y_1));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I28_un1_Y_0 (.A(
        sr_new[7]), .B(sr_prev[7]), .Y(
        SUB_13x13_medium_area_I28_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y_0 (.A(
        SUB_13x13_medium_area_I26_un1_Y_0), .B(sr_new[10]), .C(
        sr_prev[10]), .Y(SUB_13x13_medium_area_I49_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I20_S (.A(sr_new[7]), 
        .B(sr_prev[7]), .Y(N_15));
    DFN1E1C0 \deriv_out[12]  (.D(N_24), .CLK(clk_c), .CLR(n_rst_c), .E(
        deriv_enable), .Q(derivative_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I17_S (.A(sr_prev[4]), 
        .B(sr_new[4]), .Y(N_9));
    GND GND_i (.Y(GND));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I23_S (.A(sr_new[10]), 
        .B(sr_prev[10]), .Y(N_21));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I26_un1_Y_0 (.A(
        sr_new[9]), .B(sr_prev[9]), .Y(
        SUB_13x13_medium_area_I26_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I32_Y (.A(
        SUB_13x13_medium_area_I32_un1_Y_0), .B(sr_new[4]), .C(
        sr_prev[4]), .Y(N218));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I30_un1_Y_0 (.A(
        sr_new[5]), .B(sr_prev[5]), .Y(
        SUB_13x13_medium_area_I30_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y (.A(
        SUB_13x13_medium_area_I49_un1_Y_1), .B(N212), .C(
        SUB_13x13_medium_area_I49_Y_1), .Y(N204));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I32_un1_Y_0 (.A(
        sr_new[3]), .B(sr_prev[3]), .Y(
        SUB_13x13_medium_area_I32_un1_Y_0));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I31_Y (.A(sr_prev[5]), 
        .B(sr_new[5]), .C(N_13), .Y(N180));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I41_un1_Y_0 (.A(
        sr_prev[1]), .B(sr_new[1]), .C(N_5), .Y(
        SUB_13x13_medium_area_I41_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y_1 (.A(N208), .B(
        N176), .C(SUB_13x13_medium_area_I49_Y_0), .Y(
        SUB_13x13_medium_area_I49_Y_1));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I16_S (.A(sr_new[3]), 
        .B(sr_prev[3]), .Y(N_7));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y (.A(
        SUB_13x13_medium_area_I42_un1_Y_1), .B(N222), .C(
        SUB_13x13_medium_area_I42_Y_1), .Y(N212));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I27_Y (.A(sr_prev[9]), 
        .B(sr_new[9]), .C(N_21), .Y(N176));
    NOR2B un2_deriv_out_0_0_SUB_13x13_medium_area_I49_un1_Y_1 (.A(
        SUB_13x13_medium_area_I49_un1_Y_0), .B(N176), .Y(
        SUB_13x13_medium_area_I49_un1_Y_1));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I49_un1_Y_0 (.A(
        sr_new[8]), .B(sr_prev[8]), .C(N_15), .Y(
        SUB_13x13_medium_area_I49_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I41_Y (.A(
        SUB_13x13_medium_area_I41_un1_Y_0), .B(N185), .C(
        SUB_13x13_medium_area_I41_Y_0), .Y(N222));
    NOR3A un2_deriv_out_0_0_SUB_13x13_medium_area_I42_un1_Y_1 (.A(N180)
        , .B(N_9), .C(N_7), .Y(SUB_13x13_medium_area_I42_un1_Y_1));
    
endmodule


module pwm_tx_400s_32s_13s_10_1000000s_45s_1(
       off_div,
       act_ctl_5_i,
       act_ctl_5_1,
       act_ctl_5_3,
       act_ctl_5_0,
       pwm_chg_0,
       pwm_chg,
       n_rst_c,
       clk_c,
       act_ctl_5_6,
       act_ctl_5_5,
       act_ctl_5_4,
       act_ctl_5,
       primary_33_c
    );
input  [31:0] off_div;
input  act_ctl_5_i;
input  act_ctl_5_1;
input  act_ctl_5_3;
input  act_ctl_5_0;
input  pwm_chg_0;
input  pwm_chg;
input  n_rst_c;
input  clk_c;
input  act_ctl_5_6;
input  act_ctl_5_5;
input  act_ctl_5_4;
input  act_ctl_5;
output primary_33_c;

    wire N_400_0, I_140_2, I_140_1, \DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] , \DWACT_COMP0_E[1] , N_18, 
        I_20_2, \counter[7]_net_1 , N_20, I_23_3, \counter[8]_net_1 , 
        N_11, N_6, N_8, \DWACT_FDEC_E[0] , N_3, \DWACT_FDEC_E[2] , 
        N_16, N_14, \counter[6]_net_1 , N_2, \counter[2]_net_1 , 
        counter_m6_0_a2_7, counter_m6_0_a2_2, counter_m6_0_a2_1, 
        counter_m6_0_a2_6, \counter[16]_net_1 , \counter[18]_net_1 , 
        counter_m6_0_a2_4, \counter[15]_net_1 , \counter[10]_net_1 , 
        \counter[17]_net_1 , \counter[13]_net_1 , \counter[14]_net_1 , 
        \counter[11]_net_1 , \counter[12]_net_1 , counter_c18, 
        \counter[9]_net_1 , counter_c8, counter_n31, 
        \counter[31]_net_1 , counter_63_0, cur_pwm_RNI343UF1_0_net_1, 
        \counter[30]_net_1 , counter_c29, counter_n30, counter_n29, 
        \counter[29]_net_1 , counter_c28, counter_n28, counter_n28_tz, 
        \counter[27]_net_1 , counter_c26, \counter[28]_net_1 , 
        counter_n27, counter_n26, counter_n26_tz, \counter[25]_net_1 , 
        counter_c24, \counter[26]_net_1 , counter_n25, counter_n24, 
        counter_n24_tz, \counter[23]_net_1 , counter_c22, 
        \counter[24]_net_1 , counter_n23, counter_n22, counter_n22_tz, 
        \counter[21]_net_1 , counter_c20, \counter[22]_net_1 , 
        counter_n21, counter_n20, counter_n20_tz, \counter[19]_net_1 , 
        \counter[20]_net_1 , counter_n19, counter_n18, counter_c17, 
        counter_n17, counter_c16, counter_n16, counter_c15, 
        counter_n15, counter_c14, counter_n14, counter_c13, 
        counter_n13, counter_c12, counter_n12, counter_c11, 
        counter_n11, counter_c10, counter_n10, counter_n10_tz, 
        counter_n9, counter_n8, counter_n8_tz, counter_c6, counter_n7, 
        counter_n6, counter_n6_tz, \counter[5]_net_1 , counter_c4, 
        counter_n5, counter_n4, counter_n4_tz, \counter[3]_net_1 , 
        counter_c2, \counter[4]_net_1 , counter_n3, counter_n2, 
        counter_n2_tz, \counter[1]_net_1 , \counter[0]_net_1 , 
        \off_time[1] , \off_reg[1]_net_1 , \off_time[2] , 
        \off_reg[2]_net_1 , \off_time[3] , \off_reg[3]_net_1 , 
        \off_time[5] , \off_reg[5]_net_1 , \off_time[8] , 
        \off_reg[8]_net_1 , \off_time[10] , \off_reg[10]_net_1 , 
        \off_time[11] , \off_reg[11]_net_1 , \off_time[12] , 
        \off_reg[12]_net_1 , \off_time[13] , \off_reg[13]_net_1 , 
        \off_time[17] , \off_reg[17]_net_1 , \off_time[25] , 
        \off_reg[25]_net_1 , \off_time[26] , \off_reg[26]_net_1 , 
        \off_time[28] , \off_reg[28]_net_1 , \off_time[20] , 
        \off_reg[20]_net_1 , \off_time[7] , \off_reg[7]_net_1 , 
        \off_time[6] , \off_reg[6]_net_1 , \off_time[24] , 
        \off_reg[24]_net_1 , \off_time[23] , \off_reg[23]_net_1 , 
        \off_time[30] , \off_reg[30]_net_1 , \off_time[31] , 
        \off_reg[31]_net_1 , \off_time[27] , \off_reg[27]_net_1 , 
        \off_time[16] , \off_reg[16]_net_1 , \off_time[15] , 
        \off_reg[15]_net_1 , \off_time[29] , \off_reg[29]_net_1 , 
        \off_time[18] , \off_reg[18]_net_1 , \off_time[14] , 
        \off_reg[14]_net_1 , \off_time[19] , \off_reg[19]_net_1 , 
        \off_time[22] , \off_reg[22]_net_1 , \off_time[21] , 
        \off_reg[21]_net_1 , \off_time[9] , \off_reg[9]_net_1 , 
        \off_time[4] , \off_reg[4]_net_1 , \off_time[0] , 
        \off_reg[0]_net_1 , counter_n1, \counter_RNO_0[0] , 
        cur_pwm_RNO_0, \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] , N_4, N_21, N_17, N_13, 
        I_14_2, \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] , \DWACT_BL_EQUAL_0_E[3] , 
        \DWACT_BL_EQUAL_0_E[2] , \DWACT_BL_EQUAL_0_E[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] , \DWACT_COMP0_E_0[1] , 
        \DWACT_COMP0_E_0[2] , \DWACT_COMP0_E[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] , N_11_0, N_10, N_9, N_6_0, 
        N_8_0, N_7, N_5, N_2_0, N_3_0, N_4_0, N_21_0, N_20_0, N_19, 
        N_16_0, N_18_0, N_17_0, N_15, N_12, N_13_0, N_14_0, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] , 
        \DWACT_BL_EQUAL_0_E[4] , \DWACT_BL_EQUAL_0_E_0[3] , 
        \DWACT_BL_EQUAL_0_E_0[0] , \DWACT_BL_EQUAL_0_E[1] , 
        \DWACT_BL_EQUAL_0_E_0[2] , \DWACT_CMPLE_PO0_DWACT_COMP0_E[1] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[0] , N_31, N_30, N_29, N_26, 
        N_28, N_27, N_25, N_22, N_23, N_24, \ACT_LT4_E[3] , 
        \ACT_LT4_E[6] , \ACT_LT4_E[10] , \ACT_LT4_E[7] , 
        \ACT_LT4_E[8] , \ACT_LT4_E[5] , \ACT_LT4_E[4] , \ACT_LT4_E[0] , 
        \ACT_LT4_E[1] , \ACT_LT4_E[2] , \DWACT_BL_EQUAL_0_E_1[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] , 
        \DWACT_BL_EQUAL_0_E_1[0] , \DWACT_BL_EQUAL_0_E_0[1] , 
        \DWACT_BL_EQUAL_0_E_1[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] , 
        \DWACT_BL_EQUAL_0_E_2[0] , \DWACT_BL_EQUAL_0_E_1[1] , 
        \DWACT_BL_EQUAL_0_E_2[2] , \DWACT_BL_EQUAL_0_E_2[3] , 
        \DWACT_BL_EQUAL_0_E_0[4] , \DWACT_BL_EQUAL_0_E[5] , 
        \DWACT_BL_EQUAL_0_E[6] , \DWACT_BL_EQUAL_0_E[7] , 
        \DWACT_BL_EQUAL_0_E[8] , \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] , N_41, N_40, N_39, N_36, 
        N_38, N_37, N_35, N_32, N_33, N_34, \ACT_LT3_E[3] , 
        \ACT_LT3_E[4] , \ACT_LT3_E[5] , \ACT_LT3_E[0] , \ACT_LT3_E[1] , 
        \ACT_LT3_E[2] , \DWACT_BL_EQUAL_0_E_3[2] , 
        \DWACT_BL_EQUAL_0_E_2[1] , \DWACT_BL_EQUAL_0_E_3[0] , N_51, 
        N_50, N_49, N_46, N_48, N_47, N_45, N_42, N_43, N_44, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] , 
        \DWACT_BL_EQUAL_0_E_1[4] , \DWACT_BL_EQUAL_0_E_3[3] , 
        \DWACT_BL_EQUAL_0_E_4[0] , \DWACT_BL_EQUAL_0_E_3[1] , 
        \DWACT_BL_EQUAL_0_E_4[2] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] , 
        \DWACT_BL_EQUAL_0_E[12] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] , 
        \DWACT_BL_EQUAL_0_E_5[0] , \DWACT_BL_EQUAL_0_E_4[1] , 
        \DWACT_BL_EQUAL_0_E_5[2] , \DWACT_BL_EQUAL_0_E_4[3] , 
        \DWACT_BL_EQUAL_0_E_2[4] , \DWACT_BL_EQUAL_0_E_0[5] , 
        \DWACT_BL_EQUAL_0_E_0[6] , \DWACT_BL_EQUAL_0_E_0[7] , 
        \DWACT_BL_EQUAL_0_E_0[8] , \DWACT_BL_EQUAL_0_E[9] , 
        \DWACT_BL_EQUAL_0_E[10] , \DWACT_BL_EQUAL_0_E[11] , N_2_1, 
        N_5_0, GND, VCC;
    
    DFN1C0 \counter[19]  (.D(counter_n19), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[19]_net_1 ));
    AND3 un1_counter_0_I_78 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] ));
    NOR2B \counter_RNIET7L[16]  (.A(counter_c15), .B(
        \counter[16]_net_1 ), .Y(counter_c16));
    NOR3 un1_counter_2_0_I_17 (.A(\counter[20]_net_1 ), .B(
        \counter[19]_net_1 ), .C(\counter[21]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] ));
    XOR2 un1_act_ctl_I_23 (.A(act_ctl_5), .B(N_2_1), .Y(I_23_3));
    AND2A un1_counter_0_I_51 (.A(\off_time[26] ), .B(
        \counter[26]_net_1 ), .Y(\ACT_LT3_E[5] ));
    DFN1E1C0 \off_reg[28]  (.D(off_div[28]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[28]_net_1 ));
    AX1C \counter_RNO_0[2]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .C(\counter[2]_net_1 ), .Y(counter_n2_tz));
    DFN1C0 \counter[28]  (.D(counter_n28), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[28]_net_1 ));
    XNOR2 un1_counter_0_I_73 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .Y(\DWACT_BL_EQUAL_0_E_2[2] ));
    OA1A un1_counter_0_I_136 (.A(N_6_0), .B(N_8_0), .C(N_7), .Y(N_11_0)
        );
    NOR3C \counter_RNILTP7[10]  (.A(\counter[9]_net_1 ), .B(counter_c8)
        , .C(\counter[10]_net_1 ), .Y(counter_c10));
    OA1A un1_counter_0_I_132 (.A(\counter[3]_net_1 ), .B(\off_time[3] )
        , .C(N_3_0), .Y(N_7));
    DFN1E1C0 \off_reg[15]  (.D(off_div[15]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[15]_net_1 ));
    DFN1E1C0 \off_reg[26]  (.D(off_div[26]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[26]_net_1 ));
    AND3 un1_counter_0_I_14 (.A(\DWACT_BL_EQUAL_0_E[9] ), .B(
        \DWACT_BL_EQUAL_0_E[10] ), .C(\DWACT_BL_EQUAL_0_E[11] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] ));
    XA1B \counter_RNO[11]  (.A(\counter[11]_net_1 ), .B(counter_c10), 
        .C(N_400_0), .Y(counter_n11));
    DFN1C0 \counter[29]  (.D(counter_n29), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[29]_net_1 ));
    DFN1E1C0 \off_reg[5]  (.D(off_div[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[5]_net_1 ));
    NOR3 un1_counter_2_0_I_77 (.A(\counter[12]_net_1 ), .B(
        \counter[10]_net_1 ), .C(\counter[11]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] ));
    XNOR2 un1_counter_0_I_82 (.A(\counter[15]_net_1 ), .B(
        \off_time[15] ), .Y(\DWACT_BL_EQUAL_0_E_1[0] ));
    DFN1C0 \counter[11]  (.D(counter_n11), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[11]_net_1 ));
    XNOR2 un1_counter_0_I_109 (.A(\counter[6]_net_1 ), .B(
        \off_time[6] ), .Y(\DWACT_BL_EQUAL_0_E[1] ));
    NOR3C \counter_RNII5L1[2]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .C(\counter[2]_net_1 ), .Y(counter_c2));
    NOR2A un1_counter_2_0_I_118 (.A(I_14_2), .B(\counter[5]_net_1 ), 
        .Y(N_14));
    OR2A un1_counter_0_I_103 (.A(\counter[14]_net_1 ), .B(
        \off_time[14] ), .Y(N_29));
    NOR2A \counter_RNO[28]  (.A(counter_n28_tz), .B(
        cur_pwm_RNI343UF1_0_net_1), .Y(counter_n28));
    XA1B \counter_RNO[15]  (.A(\counter[15]_net_1 ), .B(counter_c14), 
        .C(N_400_0), .Y(counter_n15));
    XNOR2 un1_counter_0_I_25 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .Y(\DWACT_BL_EQUAL_0_E_3[3] ));
    AND2 un1_counter_0_I_114 (.A(\DWACT_BL_EQUAL_0_E[4] ), .B(
        \DWACT_BL_EQUAL_0_E_0[3] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] ));
    XNOR2 un1_counter_0_I_11 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .Y(\DWACT_BL_EQUAL_0_E_4[3] ));
    OR3A un1_act_ctl_I_22 (.A(act_ctl_5_1), .B(\DWACT_FDEC_E[2] ), .C(
        \DWACT_FDEC_E[0] ), .Y(N_2_1));
    OR2 \off_reg_RNIBSH9[9]  (.A(\off_reg[9]_net_1 ), .B(act_ctl_5_5), 
        .Y(\off_time[9] ));
    AX1C \counter_RNO_0[22]  (.A(\counter[21]_net_1 ), .B(counter_c20), 
        .C(\counter[22]_net_1 ), .Y(counter_n22_tz));
    XA1B \counter_RNO[7]  (.A(\counter[7]_net_1 ), .B(counter_c6), .C(
        N_400_0), .Y(counter_n7));
    OA1A un1_counter_2_0_I_125 (.A(N_16), .B(N_18), .C(N_17), .Y(N_21));
    DFN1E1C0 \off_reg[2]  (.D(off_div[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[2]_net_1 ));
    XNOR2 un1_counter_0_I_72 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .Y(\DWACT_BL_EQUAL_0_E_2[3] ));
    OA1 un1_counter_0_I_126 (.A(N_21_0), .B(N_20_0), .C(N_19), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] ));
    DFN1C0 \counter[6]  (.D(counter_n6), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[6]_net_1 ));
    AO1C un1_counter_0_I_122 (.A(\counter[7]_net_1 ), .B(\off_time[7] )
        , .C(N_12), .Y(N_18_0));
    XA1B \counter_RNO[31]  (.A(\counter[31]_net_1 ), .B(counter_63_0), 
        .C(cur_pwm_RNI343UF1_0_net_1), .Y(counter_n31));
    DFN1C0 \counter[21]  (.D(counter_n21), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[21]_net_1 ));
    AND2 un1_counter_0_I_20 (.A(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] ), .B(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] ), .Y(
        \DWACT_COMP0_E_0[1] ));
    OR2 un1_act_ctl_I_10 (.A(act_ctl_5), .B(act_ctl_5), .Y(
        \DWACT_FDEC_E[0] ));
    NOR2A \off_reg_RNI1GE8[0]  (.A(\off_reg[0]_net_1 ), .B(act_ctl_5_4)
        , .Y(\off_time[0] ));
    DFN1C0 \counter[3]  (.D(counter_n3), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[3]_net_1 ));
    DFN1C0 \counter[2]  (.D(counter_n2), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[2]_net_1 ));
    AND3 un1_counter_0_I_45 (.A(\DWACT_BL_EQUAL_0_E_3[2] ), .B(
        \DWACT_BL_EQUAL_0_E_2[1] ), .C(\DWACT_BL_EQUAL_0_E_3[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] ));
    DFN1E1C0 \off_reg[23]  (.D(off_div[23]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[23]_net_1 ));
    NOR2A \counter_RNO[8]  (.A(counter_n8_tz), .B(
        cur_pwm_RNI343UF1_0_net_1), .Y(counter_n8));
    OA1A un1_counter_2_0_I_121 (.A(\counter[8]_net_1 ), .B(I_23_3), .C(
        N_13), .Y(N_17));
    XA1B \counter_RNO[13]  (.A(\counter[13]_net_1 ), .B(counter_c12), 
        .C(N_400_0), .Y(counter_n13));
    AO1C un1_counter_0_I_57 (.A(\off_time[20] ), .B(
        \counter[20]_net_1 ), .C(N_34), .Y(N_36));
    DFN1E1C0 \off_reg[9]  (.D(off_div[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[9]_net_1 ));
    XNOR2 un1_counter_0_I_26 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(\DWACT_BL_EQUAL_0_E_4[2] ));
    AX1C \counter_RNO_0[4]  (.A(\counter[3]_net_1 ), .B(counter_c2), 
        .C(\counter[4]_net_1 ), .Y(counter_n4_tz));
    AO1C un1_counter_0_I_35 (.A(\off_time[28] ), .B(
        \counter[28]_net_1 ), .C(N_44), .Y(N_46));
    AO1 un1_counter_0_I_65 (.A(\DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] ), 
        .B(\DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] ), .C(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] ), .Y(\DWACT_COMP0_E[0] ));
    AND2 un1_counter_0_I_84 (.A(\DWACT_BL_EQUAL_0_E_1[3] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[1] ));
    DFN1C0 cur_pwm (.D(cur_pwm_RNO_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        primary_33_c));
    XA1B \counter_RNO[12]  (.A(\counter[12]_net_1 ), .B(counter_c11), 
        .C(N_400_0), .Y(counter_n12));
    NOR2B \counter_RNII50J[15]  (.A(counter_c14), .B(
        \counter[15]_net_1 ), .Y(counter_c15));
    AOI1A un1_counter_0_I_95 (.A(\ACT_LT4_E[3] ), .B(\ACT_LT4_E[6] ), 
        .C(\ACT_LT4_E[10] ), .Y(\DWACT_CMPLE_PO0_DWACT_COMP0_E[0] ));
    OA1A un1_counter_0_I_40 (.A(N_46), .B(N_48), .C(N_47), .Y(N_51));
    XA1B \counter_RNO[1]  (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(N_400_0), .Y(counter_n1));
    DFN1C0 \counter[17]  (.D(counter_n17), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[17]_net_1 ));
    NOR2 un1_counter_2_0_I_129 (.A(\counter[0]_net_1 ), .B(act_ctl_5_3)
        , .Y(N_4));
    DFN1C0 \counter[4]  (.D(counter_n4), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[4]_net_1 ));
    AO1B un1_counter_2_0_I_131 (.A(act_ctl_5_0), .B(\counter[1]_net_1 )
        , .C(N_4), .Y(N_6));
    AND2 un1_counter_0_I_30 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] ));
    NOR3C \counter_RNIVU7U[19]  (.A(\counter[19]_net_1 ), .B(
        counter_c18), .C(\counter[20]_net_1 ), .Y(counter_c20));
    OR2A un1_counter_0_I_60 (.A(\counter[23]_net_1 ), .B(
        \off_time[23] ), .Y(N_39));
    DFN1E1C0 \off_reg[11]  (.D(off_div[11]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[11]_net_1 ));
    AND2 un1_counter_0_I_29 (.A(\DWACT_BL_EQUAL_0_E_1[4] ), .B(
        \DWACT_BL_EQUAL_0_E_3[3] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] ));
    DFN1E1C0 \off_reg[22]  (.D(off_div[22]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[22]_net_1 ));
    DFN1C0 \counter[10]  (.D(counter_n10), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[10]_net_1 ));
    NOR2A un1_counter_2_0_I_19 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] ), .B(\counter[31]_net_1 )
        , .Y(\DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] ));
    NOR2A un1_counter_0_I_46 (.A(\off_time[24] ), .B(
        \counter[24]_net_1 ), .Y(\ACT_LT3_E[0] ));
    GND GND_i (.Y(GND));
    DFN1C0 \counter[13]  (.D(counter_n13), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[13]_net_1 ));
    XNOR2 un1_counter_0_I_81 (.A(\counter[16]_net_1 ), .B(
        \off_time[16] ), .Y(\DWACT_BL_EQUAL_0_E_0[1] ));
    NOR2A un1_counter_0_I_90 (.A(\off_time[18] ), .B(
        \counter[18]_net_1 ), .Y(\ACT_LT4_E[5] ));
    XNOR2 un1_counter_0_I_74 (.A(\counter[11]_net_1 ), .B(
        \off_time[11] ), .Y(\DWACT_BL_EQUAL_0_E_1[1] ));
    NOR2B un1_counter_2_0_I_140 (.A(\DWACT_COMP0_E[2] ), .B(
        \DWACT_COMP0_E[1] ), .Y(I_140_1));
    OA1A un1_counter_0_I_36 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .C(N_43), .Y(N_47));
    NOR2A \off_reg_RNITJ09[28]  (.A(\off_reg[28]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[28] ));
    XNOR2 un1_counter_0_I_66 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\DWACT_BL_EQUAL_0_E[8] ));
    AND3 un1_counter_0_I_17 (.A(\DWACT_BL_EQUAL_0_E_5[0] ), .B(
        \DWACT_BL_EQUAL_0_E_4[1] ), .C(\DWACT_BL_EQUAL_0_E_5[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] ));
    DFN1E1C0 \off_reg[17]  (.D(off_div[17]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[17]_net_1 ));
    AX1C \counter_RNO_0[10]  (.A(\counter[9]_net_1 ), .B(counter_c8), 
        .C(\counter[10]_net_1 ), .Y(counter_n10_tz));
    NOR2A \off_reg_RNINBT7[23]  (.A(\off_reg[23]_net_1 ), .B(
        act_ctl_5_5), .Y(\off_time[23] ));
    DFN1C0 \counter[12]  (.D(counter_n12), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[12]_net_1 ));
    OR2A un1_counter_0_I_130 (.A(\off_time[4] ), .B(\counter[4]_net_1 )
        , .Y(N_5));
    NOR2A \off_reg_RNIMD19[30]  (.A(\off_reg[30]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[30] ));
    NOR2B un1_counter_2_0_I_139 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E[2] )
        , .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ), .Y(
        \DWACT_COMP0_E[2] ));
    NOR2A \off_reg_RNIM9S7[13]  (.A(\off_reg[13]_net_1 ), .B(
        act_ctl_5_5), .Y(\off_time[13] ));
    NOR2A \off_reg_RNI9QH9[7]  (.A(\off_reg[7]_net_1 ), .B(act_ctl_5_5)
        , .Y(\off_time[7] ));
    DFN1C0 \counter[27]  (.D(counter_n27), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[27]_net_1 ));
    NOR3C \counter_RNIUASB1[26]  (.A(\counter[25]_net_1 ), .B(
        counter_c24), .C(\counter[26]_net_1 ), .Y(counter_c26));
    OR2A un1_counter_0_I_96 (.A(\off_time[11] ), .B(
        \counter[11]_net_1 ), .Y(N_22));
    NOR3C \counter_RNI8J6B[18]  (.A(\counter[16]_net_1 ), .B(
        \counter[18]_net_1 ), .C(counter_m6_0_a2_4), .Y(
        counter_m6_0_a2_6));
    AOI1A un1_counter_0_I_49 (.A(\ACT_LT3_E[0] ), .B(\ACT_LT3_E[1] ), 
        .C(\ACT_LT3_E[2] ), .Y(\ACT_LT3_E[3] ));
    NOR2B \counter_RNIRUMI1[29]  (.A(counter_c28), .B(
        \counter[29]_net_1 ), .Y(counter_c29));
    AX1C \counter_RNO_0[20]  (.A(\counter[19]_net_1 ), .B(counter_c18), 
        .C(\counter[20]_net_1 ), .Y(counter_n20_tz));
    DFN1C0 \counter[20]  (.D(counter_n20), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[20]_net_1 ));
    OA1A un1_counter_0_I_101 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .C(N_23), .Y(N_27));
    DFN1E1C0 \off_reg[19]  (.D(off_div[19]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[19]_net_1 ));
    NOR3C \counter_RNI5OA71[24]  (.A(\counter[23]_net_1 ), .B(
        counter_c22), .C(\counter[24]_net_1 ), .Y(counter_c24));
    XNOR2 un1_counter_0_I_71 (.A(\counter[10]_net_1 ), .B(
        \off_time[10] ), .Y(\DWACT_BL_EQUAL_0_E_2[0] ));
    OR2A un1_counter_0_I_116 (.A(\off_time[6] ), .B(\counter[6]_net_1 )
        , .Y(N_12));
    AO1C un1_counter_0_I_39 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .C(N_45), .Y(N_50));
    XA1B \counter_RNO[17]  (.A(\counter[17]_net_1 ), .B(counter_c16), 
        .C(N_400_0), .Y(counter_n17));
    XNOR2 un1_counter_0_I_69 (.A(\counter[16]_net_1 ), .B(
        \off_time[16] ), .Y(\DWACT_BL_EQUAL_0_E[6] ));
    XNOR2 un1_counter_0_I_112 (.A(\counter[9]_net_1 ), .B(
        \off_time[9] ), .Y(\DWACT_BL_EQUAL_0_E[4] ));
    OA1A un1_counter_0_I_105 (.A(N_26), .B(N_28), .C(N_27), .Y(N_31));
    DFN1C0 \counter[23]  (.D(counter_n23), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[23]_net_1 ));
    XA1B \counter_RNO[29]  (.A(\counter[29]_net_1 ), .B(counter_c28), 
        .C(cur_pwm_RNI343UF1_0_net_1), .Y(counter_n29));
    DFN1E1C0 \off_reg[25]  (.D(off_div[25]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[25]_net_1 ));
    NOR2B \counter_RNO_0[18]  (.A(counter_c16), .B(\counter[17]_net_1 )
        , .Y(counter_c17));
    DFN1C0 \counter[22]  (.D(counter_n22), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[22]_net_1 ));
    DFN1C0 \counter[15]  (.D(counter_n15), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[15]_net_1 ));
    AO1 un1_counter_0_I_107 (.A(\DWACT_CMPLE_PO0_DWACT_COMP0_E[1] ), 
        .B(\DWACT_CMPLE_PO0_DWACT_COMP0_E[2] ), .C(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] ));
    OR2A un1_counter_0_I_99 (.A(\off_time[14] ), .B(
        \counter[14]_net_1 ), .Y(N_25));
    NOR2A un1_counter_2_0_I_122 (.A(I_20_2), .B(\counter[7]_net_1 ), 
        .Y(N_18));
    AND2 un1_counter_2_0_I_115 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] ));
    XNOR2 un1_counter_0_I_108 (.A(\counter[5]_net_1 ), .B(
        \off_time[5] ), .Y(\DWACT_BL_EQUAL_0_E_0[0] ));
    AX1C \counter_RNO_0[8]  (.A(\counter[7]_net_1 ), .B(counter_c6), 
        .C(\counter[8]_net_1 ), .Y(counter_n8_tz));
    AX1C \counter_RNO_0[28]  (.A(\counter[27]_net_1 ), .B(counter_c26), 
        .C(\counter[28]_net_1 ), .Y(counter_n28_tz));
    VCC VCC_i (.Y(VCC));
    AO1C un1_counter_0_I_120 (.A(\off_time[6] ), .B(\counter[6]_net_1 )
        , .C(N_14_0), .Y(N_16_0));
    DFN1E1C0 \off_reg[31]  (.D(off_div[31]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[31]_net_1 ));
    XA1B \counter_RNO[14]  (.A(\counter[14]_net_1 ), .B(counter_c13), 
        .C(N_400_0), .Y(counter_n14));
    XNOR2 un1_counter_2_0_I_111 (.A(\counter[7]_net_1 ), .B(I_20_2), 
        .Y(\DWACT_BL_EQUAL_0_E[2] ));
    OR2 \off_reg_RNI8PH9[6]  (.A(\off_reg[6]_net_1 ), .B(act_ctl_5_5), 
        .Y(\off_time[6] ));
    DFN1E1C0 \off_reg[7]  (.D(off_div[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[7]_net_1 ));
    DFN1C0 \counter[1]  (.D(counter_n1), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[1]_net_1 ));
    XNOR2 un1_counter_0_I_2 (.A(\counter[19]_net_1 ), .B(
        \off_time[19] ), .Y(\DWACT_BL_EQUAL_0_E_5[0] ));
    MX2C cur_pwm_RNI343UF1_0 (.A(I_140_2), .B(I_140_1), .S(
        primary_33_c), .Y(cur_pwm_RNI343UF1_0_net_1));
    NOR2A \counter_RNO[26]  (.A(counter_n26_tz), .B(
        cur_pwm_RNI343UF1_0_net_1), .Y(counter_n26));
    NOR2A un1_counter_0_I_55 (.A(\off_time[19] ), .B(
        \counter[19]_net_1 ), .Y(N_34));
    AO1 un1_counter_0_I_139 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] ), .Y(\DWACT_COMP0_E_0[2] )
        );
    XA1B \counter_RNO[5]  (.A(\counter[5]_net_1 ), .B(counter_c4), .C(
        N_400_0), .Y(counter_n5));
    AO1C un1_counter_0_I_133 (.A(\counter[2]_net_1 ), .B(\off_time[2] )
        , .C(N_2_0), .Y(N_8_0));
    OR2 \off_reg_RNINAS7[14]  (.A(\off_reg[14]_net_1 ), .B(act_ctl_5_5)
        , .Y(\off_time[14] ));
    DFN1C0 \counter[25]  (.D(counter_n25), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[25]_net_1 ));
    AND2A un1_counter_0_I_87 (.A(\off_time[16] ), .B(
        \counter[16]_net_1 ), .Y(\ACT_LT4_E[2] ));
    XA1B \counter_RNO[3]  (.A(\counter[3]_net_1 ), .B(counter_c2), .C(
        N_400_0), .Y(counter_n3));
    NOR2A \off_reg_RNIRH09[26]  (.A(\off_reg[26]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[26] ));
    DFN1E1C0 \off_reg[6]  (.D(off_div[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[6]_net_1 ));
    AND3 un1_counter_0_I_28 (.A(\DWACT_BL_EQUAL_0_E_4[0] ), .B(
        \DWACT_BL_EQUAL_0_E_3[1] ), .C(\DWACT_BL_EQUAL_0_E_4[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] ));
    NOR2A \off_reg_RNIK8T7[20]  (.A(\off_reg[20]_net_1 ), .B(
        act_ctl_5_5), .Y(\off_time[20] ));
    OR2A un1_counter_0_I_50 (.A(\off_time[26] ), .B(
        \counter[26]_net_1 ), .Y(\ACT_LT3_E[4] ));
    DFN1C0 \counter[5]  (.D(counter_n5), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[5]_net_1 ));
    MX2A cur_pwm_RNO (.A(I_140_2), .B(I_140_1), .S(primary_33_c), .Y(
        cur_pwm_RNO_0));
    NOR2A \off_reg_RNIJ6S7[10]  (.A(\off_reg[10]_net_1 ), .B(
        act_ctl_5_5), .Y(\off_time[10] ));
    XNOR2 un1_counter_0_I_4 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(\DWACT_BL_EQUAL_0_E[10] ));
    XNOR2 un1_counter_0_I_23 (.A(\counter[27]_net_1 ), .B(
        \off_time[27] ), .Y(\DWACT_BL_EQUAL_0_E_4[0] ));
    NOR2A \counter_RNO[10]  (.A(counter_n10_tz), .B(
        cur_pwm_RNI343UF1_0_net_1), .Y(counter_n10));
    AND3 un1_counter_0_I_77 (.A(\DWACT_BL_EQUAL_0_E_2[0] ), .B(
        \DWACT_BL_EQUAL_0_E_1[1] ), .C(\DWACT_BL_EQUAL_0_E_2[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] ));
    XNOR2 un1_counter_0_I_3 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .Y(\DWACT_BL_EQUAL_0_E[11] ));
    XA1B \counter_RNO[21]  (.A(\counter[21]_net_1 ), .B(counter_c20), 
        .C(N_400_0), .Y(counter_n21));
    NOR2B \counter_RNINEOG[14]  (.A(counter_c13), .B(
        \counter[14]_net_1 ), .Y(counter_c14));
    XNOR2 un1_counter_0_I_6 (.A(\counter[20]_net_1 ), .B(
        \off_time[20] ), .Y(\DWACT_BL_EQUAL_0_E_4[1] ));
    OR2A un1_counter_0_I_56 (.A(\off_time[23] ), .B(
        \counter[23]_net_1 ), .Y(N_35));
    NOR2B \counter_RNITOGE[13]  (.A(counter_c12), .B(
        \counter[13]_net_1 ), .Y(counter_c13));
    NOR2A \off_reg_RNI4LH9[2]  (.A(\off_reg[2]_net_1 ), .B(act_ctl_5_5)
        , .Y(\off_time[2] ));
    AX1C \counter_RNO_0[24]  (.A(\counter[23]_net_1 ), .B(counter_c22), 
        .C(\counter[24]_net_1 ), .Y(counter_n24_tz));
    AND3 un1_counter_0_I_15 (.A(\DWACT_BL_EQUAL_0_E_0[6] ), .B(
        \DWACT_BL_EQUAL_0_E_0[7] ), .C(\DWACT_BL_EQUAL_0_E_0[8] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] ));
    AND2A un1_counter_0_I_48 (.A(\off_time[25] ), .B(
        \counter[25]_net_1 ), .Y(\ACT_LT3_E[2] ));
    NOR2A \off_reg_RNI5MH9[3]  (.A(\off_reg[3]_net_1 ), .B(act_ctl_5_5)
        , .Y(\off_time[3] ));
    NOR2A un1_counter_0_I_129 (.A(\off_time[0] ), .B(
        \counter[0]_net_1 ), .Y(N_4_0));
    XNOR2 un1_counter_0_I_9 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(\DWACT_BL_EQUAL_0_E[12] ));
    AO1 un1_counter_0_I_140 (.A(\DWACT_COMP0_E_0[1] ), .B(
        \DWACT_COMP0_E_0[2] ), .C(\DWACT_COMP0_E[0] ), .Y(I_140_2));
    OR2A un1_counter_0_I_123 (.A(\counter[9]_net_1 ), .B(\off_time[9] )
        , .Y(N_19));
    DFN1C0 \counter[16]  (.D(counter_n16), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[16]_net_1 ));
    OR2A un1_counter_0_I_38 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(N_49));
    XA1B \counter_RNO[25]  (.A(\counter[25]_net_1 ), .B(counter_c24), 
        .C(cur_pwm_RNI343UF1_0_net_1), .Y(counter_n25));
    XNOR2 un1_counter_0_I_68 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\DWACT_BL_EQUAL_0_E[7] ));
    NOR3C \counter_RNI9GNP[9]  (.A(\counter[9]_net_1 ), .B(counter_c8), 
        .C(counter_m6_0_a2_7), .Y(counter_c18));
    XNOR2 un1_act_ctl_I_14 (.A(N_5_0), .B(act_ctl_5), .Y(I_14_2));
    NOR2B \counter_RNO_0[31]  (.A(\counter[30]_net_1 ), .B(counter_c29)
        , .Y(counter_63_0));
    XNOR2 un1_counter_0_I_43 (.A(\counter[25]_net_1 ), .B(
        \off_time[25] ), .Y(\DWACT_BL_EQUAL_0_E_2[1] ));
    XOR2 un1_act_ctl_I_20 (.A(act_ctl_5), .B(N_3), .Y(I_20_2));
    AO1C un1_counter_0_I_59 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .C(N_32), .Y(N_38));
    DFN1E1C0 \off_reg[21]  (.D(off_div[21]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[21]_net_1 ));
    NOR3C \counter_RNIR1EG1[27]  (.A(\counter[27]_net_1 ), .B(
        counter_c26), .C(\counter[28]_net_1 ), .Y(counter_c28));
    AO1C un1_counter_0_I_104 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .C(N_25), .Y(N_30));
    OR2 un1_counter_2_0_I_127 (.A(\counter[1]_net_1 ), .B(act_ctl_5_3), 
        .Y(N_2));
    XNOR2 un1_counter_0_I_10 (.A(\counter[24]_net_1 ), .B(
        \off_time[24] ), .Y(\DWACT_BL_EQUAL_0_E_0[5] ));
    NOR2A un1_counter_0_I_98 (.A(\off_time[10] ), .B(
        \counter[10]_net_1 ), .Y(N_24));
    NOR2A un1_counter_0_I_33 (.A(\off_time[27] ), .B(
        \counter[27]_net_1 ), .Y(N_44));
    OA1 un1_counter_0_I_63 (.A(N_41), .B(N_40), .C(N_39), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] ));
    NOR2A \counter_RNO[6]  (.A(counter_n6_tz), .B(
        cur_pwm_RNI343UF1_0_net_1), .Y(counter_n6));
    XA1B \counter_RNO[30]  (.A(\counter[30]_net_1 ), .B(counter_c29), 
        .C(cur_pwm_RNI343UF1_0_net_1), .Y(counter_n30));
    NOR2A \off_reg_RNINE19[31]  (.A(\off_reg[31]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[31] ));
    XNOR2 un1_counter_0_I_110 (.A(\counter[8]_net_1 ), .B(
        \off_time[8] ), .Y(\DWACT_BL_EQUAL_0_E_0[3] ));
    DFN1E1C0 \off_reg[27]  (.D(off_div[27]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[27]_net_1 ));
    AND3 un1_counter_0_I_16 (.A(\DWACT_BL_EQUAL_0_E_4[3] ), .B(
        \DWACT_BL_EQUAL_0_E_2[4] ), .C(\DWACT_BL_EQUAL_0_E_0[5] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] ));
    NOR2B \counter_RNI449C[12]  (.A(counter_c11), .B(
        \counter[12]_net_1 ), .Y(counter_c12));
    OR2A un1_counter_0_I_93 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\ACT_LT4_E[8] ));
    DFN1E1C0 \off_reg[8]  (.D(off_div[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[8]_net_1 ));
    DFN1C0 \counter[26]  (.D(counter_n26), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[26]_net_1 ));
    XA1B \counter_RNO[23]  (.A(\counter[23]_net_1 ), .B(counter_c22), 
        .C(N_400_0), .Y(counter_n23));
    NOR2A \off_reg_RNISI09[27]  (.A(\off_reg[27]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[27] ));
    OA1C un1_counter_2_0_I_137 (.A(\counter[3]_net_1 ), .B(N_11), .C(
        \counter[4]_net_1 ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] ));
    OR2B un1_counter_2_0_I_133 (.A(N_2), .B(\counter[2]_net_1 ), .Y(
        N_8));
    OR2 un1_act_ctl_I_19 (.A(\DWACT_FDEC_E[2] ), .B(\DWACT_FDEC_E[0] ), 
        .Y(N_3));
    DFN1C0 \counter[14]  (.D(counter_n14), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[14]_net_1 ));
    DFN1E1C0 \off_reg[29]  (.D(off_div[29]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[29]_net_1 ));
    AND3 un1_counter_2_0_I_18 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] ));
    DFN1E1C0 \off_reg[1]  (.D(off_div[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[1]_net_1 ));
    NOR2A \counter_RNO[22]  (.A(counter_n22_tz), .B(
        cur_pwm_RNI343UF1_0_net_1), .Y(counter_n22));
    AO1C un1_counter_0_I_131 (.A(\off_time[1] ), .B(\counter[1]_net_1 )
        , .C(N_4_0), .Y(N_6_0));
    AND2 un1_counter_0_I_19 (.A(\DWACT_BL_EQUAL_0_E[12] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] ));
    XNOR2 un1_counter_0_I_42 (.A(\counter[26]_net_1 ), .B(
        \off_time[26] ), .Y(\DWACT_BL_EQUAL_0_E_3[2] ));
    AO1C un1_counter_0_I_135 (.A(\counter[3]_net_1 ), .B(\off_time[3] )
        , .C(N_5), .Y(N_10));
    DFN1E1C0 \off_reg[10]  (.D(off_div[10]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[10]_net_1 ));
    NOR2A un1_counter_0_I_85 (.A(\off_time[15] ), .B(
        \counter[15]_net_1 ), .Y(\ACT_LT4_E[0] ));
    DFN1C0 \counter[31]  (.D(counter_n31), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[31]_net_1 ));
    NOR2A \off_reg_RNIOCT7[24]  (.A(\off_reg[24]_net_1 ), .B(
        act_ctl_5_5), .Y(\off_time[24] ));
    OR2A un1_counter_0_I_32 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(N_43));
    OA1A un1_counter_0_I_62 (.A(N_36), .B(N_38), .C(N_37), .Y(N_41));
    NOR3C \counter_RNIHC05[8]  (.A(\counter[7]_net_1 ), .B(counter_c6), 
        .C(\counter[8]_net_1 ), .Y(counter_c8));
    OR3A un1_act_ctl_I_13 (.A(act_ctl_5_1), .B(act_ctl_5_1), .C(
        \DWACT_FDEC_E[0] ), .Y(N_5_0));
    NOR2A \off_reg_RNIK7S7[11]  (.A(\off_reg[11]_net_1 ), .B(
        act_ctl_5_5), .Y(\off_time[11] ));
    OA1 un1_counter_0_I_137 (.A(N_11_0), .B(N_10), .C(N_9), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] ));
    AO1 un1_counter_0_I_138 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] ));
    NOR2A un1_counter_0_I_92 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\ACT_LT4_E[7] ));
    DFN1C0 \counter[24]  (.D(counter_n24), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[24]_net_1 ));
    OR2A un1_counter_0_I_119 (.A(\off_time[9] ), .B(\counter[9]_net_1 )
        , .Y(N_15));
    NOR3 un1_counter_2_0_I_14 (.A(\counter[29]_net_1 ), .B(
        \counter[30]_net_1 ), .C(\counter[28]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] ));
    AND3 un1_counter_2_0_I_78 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ));
    XNOR2 un1_counter_0_I_80 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\DWACT_BL_EQUAL_0_E_1[2] ));
    XNOR2 un1_counter_0_I_5 (.A(\counter[27]_net_1 ), .B(
        \off_time[27] ), .Y(\DWACT_BL_EQUAL_0_E_0[8] ));
    AND3 un1_counter_0_I_113 (.A(\DWACT_BL_EQUAL_0_E_0[0] ), .B(
        \DWACT_BL_EQUAL_0_E[1] ), .C(\DWACT_BL_EQUAL_0_E_0[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] ));
    XNOR2 un1_counter_0_I_24 (.A(\counter[28]_net_1 ), .B(
        \off_time[28] ), .Y(\DWACT_BL_EQUAL_0_E_3[1] ));
    NOR2A \counter_RNO[4]  (.A(counter_n4_tz), .B(
        cur_pwm_RNI343UF1_0_net_1), .Y(counter_n4));
    AND3 un1_counter_0_I_75 (.A(\DWACT_BL_EQUAL_0_E[6] ), .B(
        \DWACT_BL_EQUAL_0_E[7] ), .C(\DWACT_BL_EQUAL_0_E[8] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] ));
    DFN1E1C0 \off_reg[14]  (.D(off_div[14]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[14]_net_1 ));
    NOR2A \off_reg_RNI6NH9[4]  (.A(\off_reg[4]_net_1 ), .B(act_ctl_5_5)
        , .Y(\off_time[4] ));
    NOR3C \counter_RNIG9P21[22]  (.A(\counter[21]_net_1 ), .B(
        counter_c20), .C(\counter[22]_net_1 ), .Y(counter_c22));
    OR2A un1_counter_2_0_I_120 (.A(N_14), .B(\counter[6]_net_1 ), .Y(
        N_16));
    NOR2B \counter_RNICG1A[11]  (.A(counter_c10), .B(
        \counter[11]_net_1 ), .Y(counter_c11));
    XA1B \counter_RNO[18]  (.A(\counter[18]_net_1 ), .B(counter_c17), 
        .C(N_400_0), .Y(counter_n18));
    NOR3 un1_counter_2_0_I_15 (.A(\counter[26]_net_1 ), .B(
        \counter[27]_net_1 ), .C(\counter[25]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] ));
    OR2A un1_counter_0_I_86 (.A(\off_time[16] ), .B(
        \counter[16]_net_1 ), .Y(\ACT_LT4_E[1] ));
    NOR2A un1_counter_2_0_I_124 (.A(I_23_3), .B(\counter[8]_net_1 ), 
        .Y(N_20));
    OA1A un1_counter_0_I_58 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .C(N_33), .Y(N_37));
    OA1A un1_counter_0_I_121 (.A(\counter[8]_net_1 ), .B(\off_time[8] )
        , .C(N_13_0), .Y(N_17_0));
    AND2 un1_counter_2_0_I_20 (.A(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] ), .B(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] ), .Y(
        \DWACT_COMP0_E[1] ));
    AX1C \counter_RNO_0[26]  (.A(\counter[25]_net_1 ), .B(counter_c24), 
        .C(\counter[26]_net_1 ), .Y(counter_n26_tz));
    XA1B \counter_RNO[27]  (.A(\counter[27]_net_1 ), .B(counter_c26), 
        .C(cur_pwm_RNI343UF1_0_net_1), .Y(counter_n27));
    OA1A un1_counter_0_I_125 (.A(N_16_0), .B(N_18_0), .C(N_17_0), .Y(
        N_21_0));
    NOR2A \off_reg_RNIL9T7[21]  (.A(\off_reg[21]_net_1 ), .B(
        act_ctl_5_5), .Y(\off_time[21] ));
    AX1C \counter_RNO_0[6]  (.A(\counter[5]_net_1 ), .B(counter_c4), 
        .C(\counter[6]_net_1 ), .Y(counter_n6_tz));
    XNOR2 un1_counter_0_I_70 (.A(\counter[15]_net_1 ), .B(
        \off_time[15] ), .Y(\DWACT_BL_EQUAL_0_E[5] ));
    OA1 un1_counter_0_I_106 (.A(N_31), .B(N_30), .C(N_29), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] ));
    NOR2B \counter_RNIJAF4[13]  (.A(\counter[13]_net_1 ), .B(
        \counter[14]_net_1 ), .Y(counter_m6_0_a2_2));
    NOR3C \counter_RNIA45K[11]  (.A(counter_m6_0_a2_2), .B(
        counter_m6_0_a2_1), .C(counter_m6_0_a2_6), .Y(
        counter_m6_0_a2_7));
    OR2 \off_reg_RNIRES7[18]  (.A(\off_reg[18]_net_1 ), .B(act_ctl_5_5)
        , .Y(\off_time[18] ));
    DFN1E1C0 \off_reg[18]  (.D(off_div[18]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[18]_net_1 ));
    AO1C un1_counter_0_I_102 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .C(N_22), .Y(N_28));
    OR2A un1_counter_2_0_I_117 (.A(\counter[7]_net_1 ), .B(I_20_2), .Y(
        N_13));
    NOR3B un1_counter_2_0_I_113 (.A(\DWACT_BL_EQUAL_0_E[2] ), .B(
        \DWACT_BL_EQUAL_0_E[0] ), .C(\counter[6]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ));
    XNOR2 un1_counter_0_I_44 (.A(\counter[24]_net_1 ), .B(
        \off_time[24] ), .Y(\DWACT_BL_EQUAL_0_E_3[0] ));
    OR2A un1_counter_0_I_53 (.A(\off_time[20] ), .B(
        \counter[20]_net_1 ), .Y(N_32));
    OR2A un1_counter_0_I_127 (.A(\off_time[1] ), .B(\counter[1]_net_1 )
        , .Y(N_2_0));
    OR2A un1_counter_0_I_34 (.A(\off_time[31] ), .B(
        \counter[31]_net_1 ), .Y(N_45));
    OR2A un1_counter_0_I_128 (.A(\counter[2]_net_1 ), .B(\off_time[2] )
        , .Y(N_3_0));
    OR2A un1_counter_0_I_89 (.A(\off_time[17] ), .B(
        \counter[17]_net_1 ), .Y(\ACT_LT4_E[4] ));
    AO1 un1_counter_0_I_64 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] ));
    DFN1E1C0 \off_reg[16]  (.D(off_div[16]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[16]_net_1 ));
    AND3 un1_counter_0_I_76 (.A(\DWACT_BL_EQUAL_0_E_2[3] ), .B(
        \DWACT_BL_EQUAL_0_E_0[4] ), .C(\DWACT_BL_EQUAL_0_E[5] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] ));
    XNOR2 un1_counter_0_I_1 (.A(\counter[23]_net_1 ), .B(
        \off_time[23] ), .Y(\DWACT_BL_EQUAL_0_E_2[4] ));
    DFN1E1C0 \off_reg[30]  (.D(off_div[30]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[30]_net_1 ));
    NOR3 un1_counter_2_0_I_75 (.A(\counter[17]_net_1 ), .B(
        \counter[18]_net_1 ), .C(\counter[16]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] ));
    NOR2A \counter_RNO[24]  (.A(counter_n24_tz), .B(
        cur_pwm_RNI343UF1_0_net_1), .Y(counter_n24));
    DFN1C0 \counter[7]  (.D(counter_n7), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[7]_net_1 ));
    AOI1A un1_counter_0_I_94 (.A(\ACT_LT4_E[7] ), .B(\ACT_LT4_E[8] ), 
        .C(\ACT_LT4_E[5] ), .Y(\ACT_LT4_E[10] ));
    NOR2A \off_reg_RNIL8S7[12]  (.A(\off_reg[12]_net_1 ), .B(
        act_ctl_5_5), .Y(\off_time[12] ));
    DFN1C0 \counter[30]  (.D(counter_n30), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[30]_net_1 ));
    NOR2B \counter_RNIF6F4[11]  (.A(\counter[11]_net_1 ), .B(
        \counter[12]_net_1 ), .Y(counter_m6_0_a2_1));
    OA1 un1_counter_0_I_41 (.A(N_51), .B(N_50), .C(N_49), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] ));
    AND3 un1_counter_0_I_18 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] ));
    OR2A un1_counter_0_I_31 (.A(\off_time[28] ), .B(
        \counter[28]_net_1 ), .Y(N_42));
    XNOR2 un1_counter_2_0_I_108 (.A(\counter[5]_net_1 ), .B(I_14_2), 
        .Y(\DWACT_BL_EQUAL_0_E[0] ));
    AO1C un1_counter_0_I_61 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .C(N_35), .Y(N_40));
    NOR2A \off_reg_RNIQG09[25]  (.A(\off_reg[25]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[25] ));
    NOR2 \counter_RNO[0]  (.A(\counter[0]_net_1 ), .B(
        cur_pwm_RNI343UF1_0_net_1), .Y(\counter_RNO_0[0] ));
    XNOR2 un1_counter_0_I_79 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\DWACT_BL_EQUAL_0_E_1[3] ));
    NOR2A \off_reg_RNIMAT7[22]  (.A(\off_reg[22]_net_1 ), .B(
        act_ctl_5_5), .Y(\off_time[22] ));
    DFN1E1C0 \off_reg[3]  (.D(off_div[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[3]_net_1 ));
    OR2 \off_reg_RNIPCS7[16]  (.A(\off_reg[16]_net_1 ), .B(act_ctl_5_5)
        , .Y(\off_time[16] ));
    NOR2A \off_reg_RNI2HE8[1]  (.A(\off_reg[1]_net_1 ), .B(act_ctl_5_4)
        , .Y(\off_time[1] ));
    DFN1E1C0 \off_reg[0]  (.D(off_div[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[0]_net_1 ));
    OR3 un1_act_ctl_I_18 (.A(act_ctl_5_1), .B(act_ctl_5_i), .C(
        act_ctl_5_1), .Y(\DWACT_FDEC_E[2] ));
    OA1B un1_counter_2_0_I_126 (.A(N_20), .B(N_21), .C(
        \counter[9]_net_1 ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ));
    OR2A un1_counter_0_I_134 (.A(\counter[4]_net_1 ), .B(\off_time[4] )
        , .Y(N_9));
    NOR3C \counter_RNIE1N6[10]  (.A(\counter[15]_net_1 ), .B(
        \counter[10]_net_1 ), .C(\counter[17]_net_1 ), .Y(
        counter_m6_0_a2_4));
    XNOR2 un1_counter_0_I_13 (.A(\counter[28]_net_1 ), .B(
        \off_time[28] ), .Y(\DWACT_BL_EQUAL_0_E[9] ));
    NOR3C \counter_RNI3PO2[4]  (.A(\counter[3]_net_1 ), .B(counter_c2), 
        .C(\counter[4]_net_1 ), .Y(counter_c4));
    OR2 \off_reg_RNIQDS7[17]  (.A(\off_reg[17]_net_1 ), .B(act_ctl_5_5)
        , .Y(\off_time[17] ));
    NOR2A un1_counter_0_I_91 (.A(\ACT_LT4_E[4] ), .B(\ACT_LT4_E[5] ), 
        .Y(\ACT_LT4_E[6] ));
    NOR2A \off_reg_RNIUK09[29]  (.A(\off_reg[29]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[29] ));
    AOI1A un1_counter_0_I_52 (.A(\ACT_LT3_E[3] ), .B(\ACT_LT3_E[4] ), 
        .C(\ACT_LT3_E[5] ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] ));
    MX2C cur_pwm_RNI343UF1 (.A(I_140_2), .B(I_140_1), .S(primary_33_c), 
        .Y(N_400_0));
    NOR2A \counter_RNO[20]  (.A(counter_n20_tz), .B(
        cur_pwm_RNI343UF1_0_net_1), .Y(counter_n20));
    NOR2A \off_reg_RNI7OH9[5]  (.A(\off_reg[5]_net_1 ), .B(act_ctl_5_5)
        , .Y(\off_time[5] ));
    NOR2A \off_reg_RNIOBS7[15]  (.A(\off_reg[15]_net_1 ), .B(
        act_ctl_5_5), .Y(\off_time[15] ));
    DFN1E1C0 \off_reg[13]  (.D(off_div[13]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[13]_net_1 ));
    XNOR2 un1_counter_0_I_27 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(\DWACT_BL_EQUAL_0_E_1[4] ));
    XNOR2 un1_counter_0_I_111 (.A(\counter[7]_net_1 ), .B(
        \off_time[7] ), .Y(\DWACT_BL_EQUAL_0_E_0[2] ));
    OR2A un1_counter_2_0_I_136 (.A(N_6), .B(N_8), .Y(N_11));
    OR2 \off_reg_RNISFS7[19]  (.A(\off_reg[19]_net_1 ), .B(act_ctl_5_5)
        , .Y(\off_time[19] ));
    AND2 un1_counter_0_I_115 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] ));
    DFN1E1C0 \off_reg[4]  (.D(off_div[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[4]_net_1 ));
    XNOR2 un1_counter_2_0_I_110 (.A(\counter[8]_net_1 ), .B(I_23_3), 
        .Y(\DWACT_BL_EQUAL_0_E[3] ));
    XNOR2 un1_counter_0_I_8 (.A(\counter[25]_net_1 ), .B(
        \off_time[25] ), .Y(\DWACT_BL_EQUAL_0_E_0[6] ));
    DFN1E1C0 \off_reg[20]  (.D(off_div[20]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[20]_net_1 ));
    NOR2A \counter_RNO[2]  (.A(counter_n2_tz), .B(
        cur_pwm_RNI343UF1_0_net_1), .Y(counter_n2));
    NOR3C \counter_RNIOGS3[5]  (.A(\counter[5]_net_1 ), .B(counter_c4), 
        .C(\counter[6]_net_1 ), .Y(counter_c6));
    DFN1C0 \counter[9]  (.D(counter_n9), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[9]_net_1 ));
    NOR3 un1_counter_2_0_I_16 (.A(\counter[24]_net_1 ), .B(
        \counter[23]_net_1 ), .C(\counter[22]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] ));
    NOR2A un1_counter_2_0_I_114 (.A(\DWACT_BL_EQUAL_0_E[3] ), .B(
        \counter[9]_net_1 ), .Y(\DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ));
    OR2A un1_counter_0_I_117 (.A(\counter[7]_net_1 ), .B(\off_time[7] )
        , .Y(N_13_0));
    XA1B \counter_RNO[19]  (.A(\counter[19]_net_1 ), .B(counter_c18), 
        .C(N_400_0), .Y(counter_n19));
    AO1C un1_counter_0_I_124 (.A(\counter[8]_net_1 ), .B(\off_time[8] )
        , .C(N_15), .Y(N_20_0));
    NOR2A un1_counter_0_I_118 (.A(\off_time[5] ), .B(
        \counter[5]_net_1 ), .Y(N_14_0));
    XNOR2 un1_counter_0_I_12 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .Y(\DWACT_BL_EQUAL_0_E_5[2] ));
    AO1 un1_counter_2_0_I_138 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] )
        , .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] ));
    NOR2A \off_reg_RNIARH9[8]  (.A(\off_reg[8]_net_1 ), .B(act_ctl_5_5)
        , .Y(\off_time[8] ));
    XA1B \counter_RNO[9]  (.A(\counter[9]_net_1 ), .B(counter_c8), .C(
        N_400_0), .Y(counter_n9));
    DFN1E1C0 \off_reg[12]  (.D(off_div[12]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[12]_net_1 ));
    AOI1A un1_counter_0_I_88 (.A(\ACT_LT4_E[0] ), .B(\ACT_LT4_E[1] ), 
        .C(\ACT_LT4_E[2] ), .Y(\ACT_LT4_E[3] ));
    OR2A un1_counter_0_I_47 (.A(\off_time[25] ), .B(
        \counter[25]_net_1 ), .Y(\ACT_LT3_E[1] ));
    DFN1C0 \counter[8]  (.D(counter_n8), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[8]_net_1 ));
    OR2A un1_counter_0_I_54 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .Y(N_33));
    AO1C un1_counter_0_I_37 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .C(N_42), .Y(N_48));
    XNOR2 un1_counter_0_I_7 (.A(\counter[26]_net_1 ), .B(
        \off_time[26] ), .Y(\DWACT_BL_EQUAL_0_E_0[7] ));
    XNOR2 un1_counter_0_I_67 (.A(\counter[14]_net_1 ), .B(
        \off_time[14] ), .Y(\DWACT_BL_EQUAL_0_E_0[4] ));
    DFN1C0 \counter[18]  (.D(counter_n18), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[18]_net_1 ));
    AO1C un1_counter_0_I_100 (.A(\off_time[11] ), .B(
        \counter[11]_net_1 ), .C(N_24), .Y(N_26));
    DFN1E1C0 \off_reg[24]  (.D(off_div[24]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[24]_net_1 ));
    AND3 un1_counter_0_I_83 (.A(\DWACT_BL_EQUAL_0_E_1[0] ), .B(
        \DWACT_BL_EQUAL_0_E_0[1] ), .C(\DWACT_BL_EQUAL_0_E_1[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] ));
    XA1B \counter_RNO[16]  (.A(\counter[16]_net_1 ), .B(counter_c15), 
        .C(N_400_0), .Y(counter_n16));
    DFN1C0 \counter[0]  (.D(\counter_RNO_0[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\counter[0]_net_1 ));
    NOR3 un1_counter_2_0_I_76 (.A(\counter[15]_net_1 ), .B(
        \counter[14]_net_1 ), .C(\counter[13]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] ));
    OR2A un1_counter_0_I_97 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .Y(N_23));
    
endmodule


module spi_clk_11s_1(
       sck_12_c,
       n_rst_c,
       clk_c
    );
output sck_12_c;
input  n_rst_c;
input  clk_c;

    wire N_8, \counter[1]_net_1 , \counter[0]_net_1 , N_6, 
        \counter[3]_net_1 , \DWACT_FINC_E[0] , cur_clk5_5, cur_clk5_3, 
        \counter[6]_net_1 , cur_clk5_4, cur_clk5_1, \counter[7]_net_1 , 
        \counter[8]_net_1 , \counter[4]_net_1 , \counter[5]_net_1 , 
        \counter[2]_net_1 , cur_clk_RNO_0, \counter_3[1] , I_5_0, 
        \counter_3[0] , \counter_3[3] , I_9_0, I_7_0, I_12_1, I_14_1, 
        I_17_1, I_20_1, I_23_1, N_2, \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[3] , N_3, N_4, \DWACT_FINC_E[1] , N_5, N_7, GND, 
        VCC;
    
    NOR2B un3_counter_I_6 (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(N_8));
    AND3 un3_counter_I_19 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\counter[6]_net_1 ), .Y(N_3));
    XOR2 un3_counter_I_20 (.A(N_3), .B(\counter[7]_net_1 ), .Y(I_20_1));
    DFN1C0 \counter[2]  (.D(I_7_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[2]_net_1 ));
    DFN1C0 \counter[7]  (.D(I_20_1), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[7]_net_1 ));
    AND3 un3_counter_I_13 (.A(\DWACT_FINC_E[0] ), .B(
        \counter[3]_net_1 ), .C(\counter[4]_net_1 ), .Y(N_5));
    AOI1 \counter_RNO[0]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(
        \counter[0]_net_1 ), .Y(\counter_3[0] ));
    DFN1C0 \counter[6]  (.D(I_17_1), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[6]_net_1 ));
    NOR3B \counter_RNIUFLE[6]  (.A(\counter[1]_net_1 ), .B(cur_clk5_3), 
        .C(\counter[6]_net_1 ), .Y(cur_clk5_5));
    VCC VCC_i (.Y(VCC));
    XOR2 un3_counter_I_12 (.A(N_6), .B(\counter[4]_net_1 ), .Y(I_12_1));
    DFN1C0 \counter[8]  (.D(I_23_1), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[8]_net_1 ));
    XOR2 un3_counter_I_23 (.A(N_2), .B(\counter[8]_net_1 ), .Y(I_23_1));
    AOI1B \counter_RNO[1]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(I_5_0), 
        .Y(\counter_3[1] ));
    AND3 un3_counter_I_22 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\DWACT_FINC_E[3] ), .Y(N_2));
    XOR2 un3_counter_I_7 (.A(N_8), .B(\counter[2]_net_1 ), .Y(I_7_0));
    NOR2B un3_counter_I_11 (.A(\counter[3]_net_1 ), .B(
        \DWACT_FINC_E[0] ), .Y(N_6));
    AND3 un3_counter_I_16 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[1] )
        , .C(\counter[5]_net_1 ), .Y(N_4));
    DFN1C0 \counter[4]  (.D(I_12_1), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[4]_net_1 ));
    XOR2 un3_counter_I_17 (.A(N_4), .B(\counter[6]_net_1 ), .Y(I_17_1));
    DFN1C0 \counter[5]  (.D(I_14_1), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[5]_net_1 ));
    AND3 un3_counter_I_8 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(N_7));
    GND GND_i (.Y(GND));
    AX1C cur_clk_RNO (.A(cur_clk5_4), .B(cur_clk5_5), .C(sck_12_c), .Y(
        cur_clk_RNO_0));
    AOI1B \counter_RNO[3]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(I_9_0), 
        .Y(\counter_3[3] ));
    AND2 un3_counter_I_21 (.A(\counter[6]_net_1 ), .B(
        \counter[7]_net_1 ), .Y(\DWACT_FINC_E[3] ));
    DFN1C0 \counter[1]  (.D(\counter_3[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[1]_net_1 ));
    DFN1C0 \counter[3]  (.D(\counter_3[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[3]_net_1 ));
    NOR3A \counter_RNI6OLE[8]  (.A(cur_clk5_1), .B(\counter[7]_net_1 ), 
        .C(\counter[8]_net_1 ), .Y(cur_clk5_4));
    NOR2 \counter_RNIVNA7[2]  (.A(\counter[5]_net_1 ), .B(
        \counter[2]_net_1 ), .Y(cur_clk5_1));
    NOR2A \counter_RNIVNA7[4]  (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(cur_clk5_3));
    AND2 un3_counter_I_15 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(\DWACT_FINC_E[1] ));
    XOR2 un3_counter_I_9 (.A(N_7), .B(\counter[3]_net_1 ), .Y(I_9_0));
    DFN1C0 cur_clk (.D(cur_clk_RNO_0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        sck_12_c));
    XOR2 un3_counter_I_14 (.A(N_5), .B(\counter[5]_net_1 ), .Y(I_14_1));
    XOR2 un3_counter_I_5 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .Y(I_5_0));
    AND3 un3_counter_I_10 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(
        \DWACT_FINC_E[0] ));
    DFN1C0 \counter[0]  (.D(\counter_3[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[0]_net_1 ));
    AND3 un3_counter_I_18 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .C(\counter[5]_net_1 ), .Y(
        \DWACT_FINC_E[2] ));
    
endmodule


module PID_controller_Z3_1(
       choose_0_0,
       choose,
       LED_FB_2,
       LED_FB_0,
       LED_5_0,
       LED_c_2,
       LED_c_0,
       LED_12_0,
       LED_15_0,
       LED_33_0,
       LED_33_2,
       LED_33_4,
       LED_33_5,
       LED_33_6,
       LED_33_7,
       primary_33_c,
       act_ctl_5,
       act_ctl_5_4,
       act_ctl_5_5,
       act_ctl_5_6,
       act_ctl_5_0,
       act_ctl_5_3,
       act_ctl_5_1,
       act_ctl_5_i,
       din_33_c,
       cs_i_1_i,
       sck_12_c,
       choose_n2,
       inc_constd,
       choose_n1,
       N_45,
       dec_constd,
       choose_n0,
       clk_c,
       n_rst_c
    );
input  choose_0_0;
input  [2:0] choose;
input  LED_FB_2;
input  LED_FB_0;
input  LED_5_0;
output LED_c_2;
output LED_c_0;
input  LED_12_0;
input  LED_15_0;
output LED_33_0;
output LED_33_2;
output LED_33_4;
output LED_33_5;
output LED_33_6;
output LED_33_7;
output primary_33_c;
input  act_ctl_5;
input  act_ctl_5_4;
input  act_ctl_5_5;
input  act_ctl_5_6;
input  act_ctl_5_0;
input  act_ctl_5_3;
input  act_ctl_5_1;
input  act_ctl_5_i;
input  din_33_c;
output cs_i_1_i;
output sck_12_c;
output choose_n2;
input  inc_constd;
output choose_n1;
input  N_45;
input  dec_constd;
output choose_n0;
input  clk_c;
input  n_rst_c;

    wire pwm_chg, sig_prev, sig_old_i_0, avg_done, N_46_1, pwm_rdy, 
        sig_prev_0, sig_old_i_0_0, sum_rdy, deriv_enable, calc_avg, 
        calc_int, pwm_enable, sum_enable, calc_error, avg_enable, 
        int_enable, pwm_chg_0, avg_enable_0, avg_enable_1, \cur_vd[0] , 
        \cur_vd[1] , \cur_vd[2] , \cur_vd[3] , \cur_vd[4] , 
        \cur_vd[5] , \cur_vd[6] , \cur_vd[7] , \cur_vd[8] , 
        \cur_vd[9] , \cur_vd[10] , \cur_vd[11] , \avg_new[0] , 
        \avg_new[1] , \avg_new[2] , \avg_new[3] , \avg_new[4] , 
        \avg_new[5] , \avg_new[6] , \avg_new[7] , \avg_new[8] , 
        \avg_new[9] , \avg_new[10] , \avg_new[11] , \avg_old[0] , 
        \avg_old[1] , \avg_old[2] , \avg_old[3] , \avg_old[4] , 
        \avg_old[5] , \avg_old[6] , \avg_old[7] , \avg_old[8] , 
        \avg_old[9] , \avg_old[10] , \avg_old[11] , \cur_error[0] , 
        \cur_error[1] , \cur_error[2] , \cur_error[3] , \cur_error[4] , 
        \cur_error[5] , \cur_error[6] , \cur_error[7] , \cur_error[8] , 
        \cur_error[9] , \cur_error[10] , \cur_error[11] , 
        \cur_error[12] , \LED_33_i[5] , \LED_33[1] , \LED_33[3] , 
        \average[2] , \average[3] , \average[4] , \average[5] , 
        \average[6] , \sr_old[0] , \sr_old[1] , \sr_old[2] , 
        \sr_old[3] , \sr_old[4] , \sr_old[5] , \sr_old[6] , 
        \sr_old[7] , \sr_old[8] , \sr_old[9] , \sr_old[10] , 
        \sr_old[11] , \sr_old[12] , \sr_new[0] , \sr_new[1] , 
        \sr_new[2] , \sr_new[3] , \sr_new[4] , \sr_new[5] , 
        \sr_new[6] , \sr_new[7] , \sr_new[8] , \sr_new[9] , 
        \sr_new[10] , \sr_new[11] , \sr_new[12] , \sr_prev[0] , 
        \sr_prev[1] , \sr_prev[2] , \sr_prev[3] , \sr_prev[4] , 
        \sr_prev[5] , \sr_prev[6] , \sr_prev[7] , \sr_prev[8] , 
        \sr_prev[9] , \sr_prev[10] , \sr_prev[11] , \sr_prev[12] , 
        \sr_new_0[12] , \sr_new_1[12] , \integral[6] , \integral[7] , 
        \integral[8] , \integral[9] , \integral[10] , \integral[11] , 
        \integral[12] , \integral[13] , \integral[14] , \integral[15] , 
        \integral[16] , \integral[17] , \integral[18] , \integral[19] , 
        \integral[20] , \integral[21] , \integral[22] , \integral[23] , 
        \integral[24] , \integral[25] , \integral_i[24] , 
        \integral_i[25] , \integral_0[25] , \integral_1[25] , 
        \derivative[12] , \sum[39] , \sum[14] , \sum[19] , \sum[20] , 
        \sum[22] , \sum[13] , \sum[18] , \sum[17] , \sum[21] , 
        \sum[23] , \sum[16] , \sum[15] , \sum[12] , \sum[11] , 
        \sum[6] , \sum[10] , \sum[9] , \sum[5] , \sum[8] , \sum[7] , 
        \sum[4] , \sum[2] , \sum[1] , \sum[0] , \sum[3] , \sum_0[39] , 
        \sum_1[39] , \sum_2[39] , vd_done, \off_div[0] , \off_div[1] , 
        \off_div[2] , \off_div[3] , \off_div[4] , \off_div[5] , 
        \off_div[6] , \off_div[7] , \off_div[8] , \off_div[9] , 
        \off_div[10] , \off_div[11] , \off_div[12] , \off_div[13] , 
        \off_div[14] , \off_div[15] , \off_div[16] , \off_div[17] , 
        \off_div[18] , \off_div[19] , \off_div[20] , \off_div[21] , 
        \off_div[22] , \off_div[23] , \off_div[24] , \off_div[25] , 
        \off_div[26] , \off_div[27] , \off_div[28] , \off_div[29] , 
        \off_div[30] , \off_div[31] , GND, VCC;
    
    pwm_ctl_400s_32s_13s_0_1_2_2 PWM_CTL (.sum_8(\sum[8] ), .sum_39(
        \sum[39] ), .sum_12(\sum[12] ), .sum_14(\sum[14] ), .sum_9(
        \sum[9] ), .sum_10(\sum[10] ), .sum_11(\sum[11] ), .sum_13(
        \sum[13] ), .sum_15(\sum[15] ), .sum_18(\sum[18] ), .sum_21(
        \sum[21] ), .sum_22(\sum[22] ), .sum_23(\sum[23] ), .sum_16(
        \sum[16] ), .sum_17(\sum[17] ), .sum_20(\sum[20] ), .sum_19(
        \sum[19] ), .sum_1_d0(\sum[1] ), .sum_0_d0(\sum[0] ), 
        .sum_2_d0(\sum[2] ), .sum_7(\sum[7] ), .sum_6(\sum[6] ), 
        .sum_5(\sum[5] ), .sum_4(\sum[4] ), .sum_3(\sum[3] ), .off_div({
        \off_div[31] , \off_div[30] , \off_div[29] , \off_div[28] , 
        \off_div[27] , \off_div[26] , \off_div[25] , \off_div[24] , 
        \off_div[23] , \off_div[22] , \off_div[21] , \off_div[20] , 
        \off_div[19] , \off_div[18] , \off_div[17] , \off_div[16] , 
        \off_div[15] , \off_div[14] , \off_div[13] , \off_div[12] , 
        \off_div[11] , \off_div[10] , \off_div[9] , \off_div[8] , 
        \off_div[7] , \off_div[6] , \off_div[5] , \off_div[4] , 
        \off_div[3] , \off_div[2] , \off_div[1] , \off_div[0] }), 
        .sum_2_0(\sum_2[39] ), .sum_1_0(\sum_1[39] ), .sum_0_0(
        \sum_0[39] ), .n_rst_c(n_rst_c), .clk_c(clk_c), .pwm_rdy(
        pwm_rdy), .pwm_enable(pwm_enable));
    integral_calc_13s_4_0 AVG_CALC (.avg_old({\avg_old[11] , 
        \avg_old[10] , \avg_old[9] , \avg_old[8] , \avg_old[7] , 
        \avg_old[6] , \avg_old[5] , \avg_old[4] , \avg_old[3] , 
        \avg_old[2] , \avg_old[1] , \avg_old[0] }), .avg_new({
        \avg_new[11] , \avg_new[10] , \avg_new[9] , \avg_new[8] , 
        \avg_new[7] , \avg_new[6] , \avg_new[5] , \avg_new[4] , 
        \avg_new[3] , \avg_new[2] , \avg_new[1] , \avg_new[0] }), 
        .LED_15_0(LED_15_0), .LED_12_0(LED_12_0), .LED_c_2(LED_c_2), 
        .LED_c_0(LED_c_0), .LED_5_0(LED_5_0), .LED_FB_2(LED_FB_2), 
        .LED_FB_0(LED_FB_0), .choose({choose[2], choose[1], choose[0]})
        , .choose_0_0(choose_0_0), .average({\average[6] , 
        \average[5] , \average[4] , \average[3] , \average[2] }), 
        .LED_33({LED_33_7, LED_33_6, LED_33_5, LED_33_4, \LED_33[3] , 
        LED_33_2, \LED_33[1] , LED_33_0}), .LED_33_i_0(\LED_33_i[5] ), 
        .calc_avg(calc_avg), .avg_done(avg_done), .choose_n0(choose_n0)
        , .dec_constd(dec_constd), .N_45(N_45), .choose_n1(choose_n1), 
        .inc_constd(inc_constd), .choose_n2(choose_n2), .n_rst_c(
        n_rst_c), .clk_c(clk_c));
    error_sr_13s_5s_0 AVGSR (.cur_vd({\cur_vd[11] , \cur_vd[10] , 
        \cur_vd[9] , \cur_vd[8] , \cur_vd[7] , \cur_vd[6] , 
        \cur_vd[5] , \cur_vd[4] , \cur_vd[3] , \cur_vd[2] , 
        \cur_vd[1] , \cur_vd[0] }), .avg_new({\avg_new[11] , 
        \avg_new[10] , \avg_new[9] , \avg_new[8] , \avg_new[7] , 
        \avg_new[6] , \avg_new[5] , \avg_new[4] , \avg_new[3] , 
        \avg_new[2] , \avg_new[1] , \avg_new[0] }), .avg_old({
        \avg_old[11] , \avg_old[10] , \avg_old[9] , \avg_old[8] , 
        \avg_old[7] , \avg_old[6] , \avg_old[5] , \avg_old[4] , 
        \avg_old[3] , \avg_old[2] , \avg_old[1] , \avg_old[0] }), 
        .avg_enable_1(avg_enable_1), .avg_enable_0(avg_enable_0), 
        .avg_enable(avg_enable), .n_rst_c(n_rst_c), .clk_c(clk_c));
    error_sr_13s_64s_0 INTSR (.sr_old({\sr_old[12] , \sr_old[11] , 
        \sr_old[10] , \sr_old[9] , \sr_old[8] , \sr_old[7] , 
        \sr_old[6] , \sr_old[5] , \sr_old[4] , \sr_old[3] , 
        \sr_old[2] , \sr_old[1] , \sr_old[0] }), .sr_new({\sr_new[12] , 
        \sr_new[11] , \sr_new[10] , \sr_new[9] , \sr_new[8] , 
        \sr_new[7] , \sr_new[6] , \sr_new[5] , \sr_new[4] , 
        \sr_new[3] , \sr_new[2] , \sr_new[1] , \sr_new[0] }), 
        .cur_error({\cur_error[12] , \cur_error[11] , \cur_error[10] , 
        \cur_error[9] , \cur_error[8] , \cur_error[7] , \cur_error[6] , 
        \cur_error[5] , \cur_error[4] , \cur_error[3] , \cur_error[2] , 
        \cur_error[1] , \cur_error[0] }), .sr_prev({\sr_prev[12] , 
        \sr_prev[11] , \sr_prev[10] , \sr_prev[9] , \sr_prev[8] , 
        \sr_prev[7] , \sr_prev[6] , \sr_prev[5] , \sr_prev[4] , 
        \sr_prev[3] , \sr_prev[2] , \sr_prev[1] , \sr_prev[0] }), 
        .sr_new_0_0(\sr_new_0[12] ), .sr_new_1_0(\sr_new_1[12] ), 
        .int_enable(int_enable), .n_rst_c(n_rst_c), .clk_c(clk_c));
    controller_Z1_4_0 CONTROLLER (.pwm_chg(pwm_chg), .sig_prev_0(
        sig_prev), .sig_old_i_0_0(sig_old_i_0), .avg_done(avg_done), 
        .N_46_1(N_46_1), .pwm_rdy(pwm_rdy), .sig_prev(sig_prev_0), 
        .sig_old_i_0(sig_old_i_0_0), .sum_rdy(sum_rdy), .deriv_enable(
        deriv_enable), .calc_avg(calc_avg), .calc_int(calc_int), 
        .pwm_enable(pwm_enable), .sum_enable(sum_enable), .calc_error(
        calc_error), .avg_enable(avg_enable), .int_enable(int_enable), 
        .pwm_chg_0(pwm_chg_0), .avg_enable_0(avg_enable_0), .n_rst_c(
        n_rst_c), .clk_c(clk_c), .avg_enable_1(avg_enable_1));
    sig_gen_2 FM_CYCLE (.primary_33_c(primary_33_c), .n_rst_c(n_rst_c), 
        .clk_c(clk_c), .sig_old_i_0(sig_old_i_0), .sig_prev(sig_prev));
    pid_sum_13s_4_0 SUM (.integral_i({\integral_i[25] , 
        \integral_i[24] }), .sr_new({\sr_new[12] , \sr_new[11] , 
        \sr_new[10] , \sr_new[9] , \sr_new[8] , \sr_new[7] , 
        \sr_new[6] , \sr_new[5] , \sr_new[4] , \sr_new[3] , 
        \sr_new[2] , \sr_new[1] , \sr_new[0] }), .integral({
        \integral[25] , \integral[24] , \integral[23] , \integral[22] , 
        \integral[21] , \integral[20] , \integral[19] , \integral[18] , 
        \integral[17] , \integral[16] , \integral[15] , \integral[14] , 
        \integral[13] , \integral[12] , \integral[11] , \integral[10] , 
        \integral[9] , \integral[8] , \integral[7] , \integral[6] }), 
        .derivative_0(\derivative[12] ), .sr_new_0_0(\sr_new_0[12] ), 
        .sr_new_1_0(\sr_new_1[12] ), .integral_0_0(\integral_0[25] ), 
        .integral_1_0(\integral_1[25] ), .sum_39(\sum[39] ), .sum_14(
        \sum[14] ), .sum_19(\sum[19] ), .sum_20(\sum[20] ), .sum_22(
        \sum[22] ), .sum_13(\sum[13] ), .sum_18(\sum[18] ), .sum_17(
        \sum[17] ), .sum_21(\sum[21] ), .sum_23(\sum[23] ), .sum_16(
        \sum[16] ), .sum_15(\sum[15] ), .sum_12(\sum[12] ), .sum_11(
        \sum[11] ), .sum_6(\sum[6] ), .sum_10(\sum[10] ), .sum_9(
        \sum[9] ), .sum_5(\sum[5] ), .sum_8(\sum[8] ), .sum_7(\sum[7] )
        , .sum_4(\sum[4] ), .sum_2_d0(\sum[2] ), .sum_1_d0(\sum[1] ), 
        .sum_0_d0(\sum[0] ), .sum_3(\sum[3] ), .sum_0_0(\sum_0[39] ), 
        .sum_1_0(\sum_1[39] ), .sum_2_0(\sum_2[39] ), .sum_enable(
        sum_enable), .sum_rdy(sum_rdy), .n_rst_c(n_rst_c), .clk_c(
        clk_c));
    sig_gen_1 VD_SIG (.vd_done(vd_done), .n_rst_c(n_rst_c), .clk_c(
        clk_c), .sig_old_i_0(sig_old_i_0_0), .sig_prev(sig_prev_0));
    spi_rx_12s_1 SPI (.cur_vd({\cur_vd[11] , \cur_vd[10] , \cur_vd[9] , 
        \cur_vd[8] , \cur_vd[7] , \cur_vd[6] , \cur_vd[5] , 
        \cur_vd[4] , \cur_vd[3] , \cur_vd[2] , \cur_vd[1] , 
        \cur_vd[0] }), .vd_done(vd_done), .cs_i_1_i(cs_i_1_i), 
        .sck_12_c(sck_12_c), .n_rst_c(n_rst_c), .din_33_c(din_33_c));
    integral_calc_13s_0_4_0 INTCALC (.sr_new({\sr_new[12] , 
        \sr_new[11] , \sr_new[10] , \sr_new[9] , \sr_new[8] , 
        \sr_new[7] , \sr_new[6] , \sr_new[5] , \sr_new[4] , 
        \sr_new[3] , \sr_new[2] , \sr_new[1] , \sr_new[0] }), .sr_old({
        \sr_old[12] , \sr_old[11] , \sr_old[10] , \sr_old[9] , 
        \sr_old[8] , \sr_old[7] , \sr_old[6] , \sr_old[5] , 
        \sr_old[4] , \sr_old[3] , \sr_old[2] , \sr_old[1] , 
        \sr_old[0] }), .sr_new_1_0(\sr_new_1[12] ), .sr_new_0_0(
        \sr_new_0[12] ), .integral({\integral[25] , \integral[24] , 
        \integral[23] , \integral[22] , \integral[21] , \integral[20] , 
        \integral[19] , \integral[18] , \integral[17] , \integral[16] , 
        \integral[15] , \integral[14] , \integral[13] , \integral[12] , 
        \integral[11] , \integral[10] , \integral[9] , \integral[8] , 
        \integral[7] , \integral[6] }), .integral_i({\integral_i[25] , 
        \integral_i[24] }), .integral_0_0(\integral_0[25] ), 
        .integral_1_0(\integral_1[25] ), .calc_int(calc_int), .N_46_1(
        N_46_1), .n_rst_c(n_rst_c), .clk_c(clk_c));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    error_calc_13s_12s_4_0 EC (.cur_error({\cur_error[12] , 
        \cur_error[11] , \cur_error[10] , \cur_error[9] , 
        \cur_error[8] , \cur_error[7] , \cur_error[6] , \cur_error[5] , 
        \cur_error[4] , \cur_error[3] , \cur_error[2] , \cur_error[1] , 
        \cur_error[0] }), .LED_33_i_0(\LED_33_i[5] ), .LED_33({
        LED_33_7, LED_33_6, LED_33_5, LED_33_4, \LED_33[3] , LED_33_2, 
        \LED_33[1] , LED_33_0}), .average({\average[6] , \average[5] , 
        \average[4] , \average[3] , \average[2] }), .calc_error(
        calc_error), .n_rst_c(n_rst_c), .clk_c(clk_c));
    derivative_calc_13s_4_0 DCALC (.derivative_0(\derivative[12] ), 
        .sr_prev({\sr_prev[12] , \sr_prev[11] , \sr_prev[10] , 
        \sr_prev[9] , \sr_prev[8] , \sr_prev[7] , \sr_prev[6] , 
        \sr_prev[5] , \sr_prev[4] , \sr_prev[3] , \sr_prev[2] , 
        \sr_prev[1] , \sr_prev[0] }), .sr_new({\sr_new[11] , 
        \sr_new[10] , \sr_new[9] , \sr_new[8] , \sr_new[7] , 
        \sr_new[6] , \sr_new[5] , \sr_new[4] , \sr_new[3] , 
        \sr_new[2] , \sr_new[1] , \sr_new[0] }), .sr_new_1_0(
        \sr_new_1[12] ), .deriv_enable(deriv_enable), .n_rst_c(n_rst_c)
        , .clk_c(clk_c));
    pwm_tx_400s_32s_13s_10_1000000s_45s_1 PWM_TX (.off_div({
        \off_div[31] , \off_div[30] , \off_div[29] , \off_div[28] , 
        \off_div[27] , \off_div[26] , \off_div[25] , \off_div[24] , 
        \off_div[23] , \off_div[22] , \off_div[21] , \off_div[20] , 
        \off_div[19] , \off_div[18] , \off_div[17] , \off_div[16] , 
        \off_div[15] , \off_div[14] , \off_div[13] , \off_div[12] , 
        \off_div[11] , \off_div[10] , \off_div[9] , \off_div[8] , 
        \off_div[7] , \off_div[6] , \off_div[5] , \off_div[4] , 
        \off_div[3] , \off_div[2] , \off_div[1] , \off_div[0] }), 
        .act_ctl_5_i(act_ctl_5_i), .act_ctl_5_1(act_ctl_5_1), 
        .act_ctl_5_3(act_ctl_5_3), .act_ctl_5_0(act_ctl_5_0), 
        .pwm_chg_0(pwm_chg_0), .pwm_chg(pwm_chg), .n_rst_c(n_rst_c), 
        .clk_c(clk_c), .act_ctl_5_6(act_ctl_5_6), .act_ctl_5_5(
        act_ctl_5_5), .act_ctl_5_4(act_ctl_5_4), .act_ctl_5(act_ctl_5), 
        .primary_33_c(primary_33_c));
    spi_clk_11s_1 SPICLK (.sck_12_c(sck_12_c), .n_rst_c(n_rst_c), 
        .clk_c(clk_c));
    
endmodule


module pwm_ctl_400s_32s_13s_0_1_2_4(
       sum_8,
       sum_39,
       sum_10,
       sum_11,
       sum_12,
       sum_13,
       sum_14,
       sum_16,
       sum_17,
       sum_18,
       sum_19,
       sum_20,
       sum_21,
       sum_22,
       sum_23,
       sum_15,
       sum_9,
       sum_0_d0,
       sum_2_d0,
       sum_1_d0,
       sum_7,
       sum_6,
       sum_4,
       sum_3,
       sum_5,
       LED_33_0,
       LED_33_2,
       LED_33_5,
       LED_FB_0,
       LED_FB_2,
       LED_FB_5,
       LED_5_0,
       LED_5_2,
       LED_5_3,
       LED_5_5,
       choose,
       LED_c_0,
       LED_c_2,
       LED_c_5,
       LED_15_0,
       LED_15_2,
       LED_15_3,
       LED_15_5,
       LED_12_0,
       LED_12_2,
       LED_12_3,
       LED_12_5,
       choose_0_0,
       off_div,
       sum_1_0,
       sum_0_0,
       sum_2_0,
       state,
       n_rst_c,
       clk_c,
       N_45,
       pwm_enable
    );
input  sum_8;
input  sum_39;
input  sum_10;
input  sum_11;
input  sum_12;
input  sum_13;
input  sum_14;
input  sum_16;
input  sum_17;
input  sum_18;
input  sum_19;
input  sum_20;
input  sum_21;
input  sum_22;
input  sum_23;
input  sum_15;
input  sum_9;
input  sum_0_d0;
input  sum_2_d0;
input  sum_1_d0;
input  sum_7;
input  sum_6;
input  sum_4;
input  sum_3;
input  sum_5;
input  LED_33_0;
input  LED_33_2;
input  LED_33_5;
input  LED_FB_0;
input  LED_FB_2;
input  LED_FB_5;
input  LED_5_0;
input  LED_5_2;
input  LED_5_3;
input  LED_5_5;
input  [2:0] choose;
output LED_c_0;
output LED_c_2;
output LED_c_5;
input  LED_15_0;
input  LED_15_2;
input  LED_15_3;
input  LED_15_5;
input  LED_12_0;
input  LED_12_2;
input  LED_12_3;
input  LED_12_5;
input  choose_0_0;
output [31:0] off_div;
input  sum_1_0;
input  sum_0_0;
input  sum_2_0;
output [1:0] state;
input  n_rst_c;
input  clk_c;
output N_45;
input  pwm_enable;

    wire \state_d_0[2] , un1_state_2_0, un5lt31, 
        next_off_div_2_sqmuxa_10, N_16, \DWACT_FINC_E[4] , N_13, 
        \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , ADD_32x32_fast_I321_Y_0, 
        ADD_32x32_fast_I258_Y_0_1, ADD_32x32_fast_I258_Y_0_0, N482, 
        ADD_32x32_fast_I317_Y_0, ADD_32x32_fast_I258_Y_0_a5_1, 
        ADD_32x32_fast_I258_Y_0_a5_0, N483, 
        ADD_32x32_fast_I258_Y_0_o5_0, N490, N486, 
        ADD_32x32_fast_I313_Y_0, ADD_32x32_fast_I258_Y_0_a3_0, N491, 
        N487, ADD_32x32_fast_I320_Y_0, ADD_32x32_fast_I258_Y_0_o3_1, 
        N560, N567, ADD_32x32_fast_I258_Y_0_o3_0, N494, N498, 
        ADD_32x32_fast_I259_Y_3, N612, N627, ADD_32x32_fast_I259_Y_2, 
        N484, ADD_32x32_fast_I259_Y_0, N553, ADD_32x32_fast_I318_Y_0, 
        ADD_32x32_fast_I319_Y_0, ADD_32x32_fast_I258_Y_0_a3_0_0, N568, 
        ADD_32x32_fast_I316_Y_0, ADD_32x32_fast_I314_Y_0, 
        ADD_32x32_fast_I315_Y_0, ADD_32x32_fast_I261_Y_2, N616, N631, 
        ADD_32x32_fast_I261_Y_1, N488, N557, ADD_32x32_fast_I260_Y_2, 
        N614, N629, ADD_32x32_fast_I260_Y_1, N555, 
        ADD_32x32_fast_I312_Y_0, ADD_32x32_fast_I304_Y_0, 
        \sum_adj[22]_net_1 , ADD_32x32_fast_I259_un1_Y_0, N628, 
        ADD_32x32_fast_I242_Y_0, N583, N576, N575, 
        ADD_32x32_fast_I311_Y_0, ADD_32x32_fast_I310_Y_0, 
        ADD_32x32_fast_I309_Y_0, ADD_32x32_fast_I263_Y_1, N620, N635, 
        ADD_32x32_fast_I263_Y_0, N561, ADD_32x32_fast_I265_Y_0, N565, 
        ADD_32x32_fast_I264_Y_1, N622, N637, ADD_32x32_fast_I264_Y_0, 
        N563, ADD_32x32_fast_I306_Y_0, ADD_32x32_fast_I308_Y_0, 
        ADD_32x32_fast_I307_Y_0, ADD_32x32_fast_I302_Y_0, 
        \sum_adj[20]_net_1 , ADD_32x32_fast_I303_Y_0, 
        \un1_sum_adj[13] , ADD_32x32_fast_I260_un1_Y_0, N630, 
        ADD_32x32_fast_I261_un1_Y_0, N632, ADD_32x32_fast_I242_un1_Y_0, 
        N584, ADD_32x32_fast_I301_Y_0, \sum_adj[19]_net_1 , 
        ADD_32x32_fast_I269_Y_0, N647, ADD_32x32_fast_I300_Y_0, 
        \un1_sum_adj[10] , ADD_32x32_fast_I299_Y_0, \un1_sum_adj[9] , 
        ADD_32x32_fast_I298_Y_0, \un1_sum_adj[8] , 
        ADD_32x32_fast_I270_Y_1, ADD_32x32_fast_I270_un1_Y_0, N599, 
        ADD_32x32_fast_I270_Y_0, ADD_32x32_fast_I263_un1_Y_0, N636, 
        ADD_32x32_fast_I264_un1_Y_0, N638, ADD_32x32_fast_I265_un1_Y_0, 
        N582, N574, N624, ADD_32x32_fast_I296_Y_0, \un1_sum_adj[6] , 
        ADD_32x32_fast_I271_Y_0, ADD_32x32_fast_I271_un1_Y_0, 
        ADD_32x32_fast_I272_Y_0, ADD_32x32_fast_I272_un1_Y_0, 
        ADD_32x32_fast_I295_Y_0, \sum_adj[13]_net_1 , 
        ADD_32x32_fast_I294_Y_0, \un1_sum_adj[4] , 
        ADD_32x32_fast_I269_un1_Y_0, N648, ADD_32x32_fast_I293_Y_0, 
        \sum_adj[11]_net_1 , N650, N634, N538, N654, 
        ADD_32x32_fast_I273_un1_Y_0, N590, N598, \un1_sum_adj[0] , 
        N586, N594, N601, ADD_32x32_fast_I292_Y_0, \un1_sum_adj[2] , 
        next_off_div_2_sqmuxa_9, next_off_div37, 
        next_off_div_2_sqmuxa_6, next_off_div_2_sqmuxa_5, 
        next_off_div_2_sqmuxa_7, next_off_div_2_sqmuxa_4, 
        next_off_div_2_sqmuxa_2, ADD_32x32_fast_I291_Y_0, 
        \sum_adj[9]_net_1 , un5lto20_2, un5lto20_1, 
        ADD_32x32_fast_I157_Y_1, ADD_32x32_fast_I157_Y_0, N485, 
        un5lto14_2, un5lto14_1, un1_off_divlto31_22, 
        un1_off_divlto31_15, un1_off_divlto31_14, un1_off_divlto31_20, 
        un1_off_divlto31_21, un1_off_divlto31_13, un1_off_divlto31_12, 
        un1_off_divlto31_17, un1_off_divlto31_10, un1_off_divlto31_9, 
        un1_off_divlt31, un1_off_divlto31_0, un5lto9, 
        un1_off_divlto31_8, un1_off_divlto31_6, un1_off_divlto31_4, 
        un1_off_divlto31_2, un5lto7_1, N_5, N781, \un1_off_div_1[18] , 
        I236_un1_Y, \un1_off_div_1[19] , I234_un1_Y, 
        \un1_off_div_1[10] , N796, N749, N_6, N556, N753, N787, 
        I265_un1_Y, N802, N763, I224_un1_Y, N755, N790, N489, N558, 
        un1_off_div, I273_un1_Y, N779, N639, I240_un1_Y, un5lt16, 
        \un1_off_div_1[5] , N661, N759, I269_un1_Y, N663, 
        \un1_off_div_1[15] , \un1_sum_adj[15] , \un1_off_div_1[0] , 
        \un1_off_div_1[3] , \un1_off_div_1[17] , I238_un1_Y, 
        \un1_off_div_1[20] , \un1_off_div_1[7] , \un1_sum_adj[7] , 
        N657, un5lt9, un5lto4, un5lt4, N769, I230_un1_Y, I268_un1_Y, 
        N646, N767, I228_un1_Y, I267_un1_Y, N644, N659, N761, N799, 
        N751, N784, N493, \next_off_div[1] , \state_d[2] , 
        \next_off_div[2] , \next_off_div[4] , \next_off_div[6] , 
        \next_off_div[9] , \next_off_div[13] , \next_off_div[21] , 
        \next_off_div[22] , \next_off_div[25] , \next_off_div[30] , 
        N395, N401, N404, N405, N407, N408, N410, N519, N414, N520, 
        N521, N522, N523, N524, N525, N526, N398, N527, N399, N528, 
        N529, N530, N392, N517, N518, N587, N589, N593, N532, N533, 
        N643, N389, N393, N413, N417, N383, N386, N387, N390, 
        \sum_adj[10]_net_1 , N416, N419, N420, N514, N515, N516, N531, 
        N534, N535, N536, N537, \sum_adj[8]_net_1 , N511, N510, N579, 
        N580, N588, N591, N592, N595, N596, N597, I150_un1_Y, N571, 
        N564, N572, N645, N649, N653, N655, I204_un1_Y, I249_un1_Y, 
        \nsum_adj_11[10] , I_28_2, \nsum_adj_11[11] , I_32_2, 
        \nsum_adj_11[12] , I_35_2, \nsum_adj_11[13] , I_37_2, 
        \nsum_adj_11[14] , I_40_2, \nsum_adj_11[16] , I_46_2, 
        \nsum_adj_11[17] , I_49_2, \nsum_adj_11[18] , I_53_2, 
        \nsum_adj_11[19] , I_56_2, \nsum_adj_11[20] , I_59_2, 
        \nsum_adj_11[21] , I_62_2, \nsum_adj_11[22] , I_65_2, 
        \nsum_adj_11[23] , I_70_2, \sum_adj[17]_net_1 , 
        \sum_adj[16]_net_1 , \sum_adj[15]_net_1 , \sum_adj[14]_net_1 , 
        \sum_adj[12]_net_1 , N_311_i, un5lt14, \next_off_div[20] , 
        next_off_div_1_sqmuxa, \next_off_div[17] , \next_off_div[7] , 
        \next_off_div[3] , next_off_div_0_sqmuxa, \next_off_div[0] , 
        \state_ns[0] , state_176_d, N_97, N_99, N_100, N_102, N_42, 
        N_34, N_44, N_36, N_37, N_47, N_39, N_66, N_50, N_58, N_68, 
        N_52, N_60, N_71, N_55, N_63, \next_off_div[15] , 
        \sum_adj[21]_net_1 , \sum_adj[23]_net_1 , N581, N573, N566, 
        N426, N422, N425, N509, N429, N508, N428, N513, N512, 
        \next_off_div[14] , \next_off_div[26] , \next_off_div[12] , 
        un1_state_2, \next_off_div[5] , N507, N432, N506, 
        \next_off_div[16] , \nsum_adj_11[15] , I_43_2, 
        \next_off_div[28] , N492, N496, N497, \next_off_div[31] , 
        \next_off_div[29] , \next_off_div[24] , \next_off_div[23] , 
        \next_off_div[8] , \nsum_adj_11[9] , I_26_2, \nsum_adj_11[8] , 
        I_23_8, N505, N502, N499, N503, N562, N570, N577, N569, N504, 
        N501, N500, N495, \next_off_div[10] , \next_off_div[18] , 
        \next_off_div[19] , \sum_adj[18]_net_1 , N793, I247_un1_Y, 
        N651, I196_un1_Y, N585, N578, \next_off_div[27] , 
        \next_off_div[11] , N_2, \DWACT_FINC_E[29] , 
        \DWACT_FINC_E[13] , \DWACT_FINC_E[33] , \DWACT_FINC_E[34] , 
        \DWACT_FINC_E[2] , \DWACT_FINC_E[5] , \DWACT_FINC_E[15] , N_3, 
        \DWACT_FINC_E[28] , \DWACT_FINC_E[16] , N_4, N_5_0, 
        \DWACT_FINC_E[14] , N_6_0, \DWACT_FINC_E[9] , 
        \DWACT_FINC_E[12] , N_7, \DWACT_FINC_E[10] , \DWACT_FINC_E[0] , 
        N_8, \DWACT_FINC_E[11] , N_9, N_10, N_11, \DWACT_FINC_E[8] , 
        N_12, N_14, N_15, \DWACT_FINC_E[3] , N_17, GND, VCC;
    
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I59_Y (.A(sum_1_0), .B(
        off_div[17]), .C(N432), .Y(N505));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I10_P0N (.A(\un1_sum_adj[10] )
        , .B(off_div[10]), .Y(N414));
    NOR2A \LED_2[2]  (.A(LED_5_2), .B(choose[2]), .Y(N_36));
    DFN1C0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(state[0]));
    DFN1E0C0 \off_div[29]  (.D(\next_off_div[29] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[29]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y_0 (.A(N555), .B(N563), 
        .Y(ADD_32x32_fast_I264_Y_0));
    DFN1E0C0 \off_div[26]  (.D(\next_off_div[26] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[26]));
    NOR3A \off_div_RNIDHI11[24]  (.A(state[0]), .B(off_div[24]), .C(
        off_div[29]), .Y(next_off_div_2_sqmuxa_5));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I247_Y (.A(I247_un1_Y), .B(
        N651), .Y(N796));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I108_Y (.A(N496), .B(N492), 
        .Y(N557));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I47_Y (.A(off_div[23]), .B(
        off_div[22]), .C(sum_1_0), .Y(N493));
    NOR2A \state_RNIPD9M[0]  (.A(state[1]), .B(state[0]), .Y(
        \state_d_0[2] ));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I3_P0N (.A(sum_0_0), .B(
        \sum_adj[11]_net_1 ), .C(off_div[3]), .Y(N393));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I165_Y (.A(N489), .B(N493), 
        .C(N562), .Y(N620));
    XNOR2 un13_nsum_adj_I_49 (.A(sum_17), .B(N_8), .Y(I_49_2));
    NOR3 un13_nsum_adj_I_10 (.A(sum_0_d0), .B(sum_2_d0), .C(sum_1_d0), 
        .Y(\DWACT_FINC_E[0] ));
    DFN1E0C0 \off_div[31]  (.D(\next_off_div[31] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[31]));
    MX2 \LED_6[2]  (.A(N_52), .B(N_60), .S(choose[1]), .Y(N_68));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I149_Y (.A(N537), .B(N533), 
        .Y(N598));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I135_Y (.A(N523), .B(N519), 
        .Y(N584));
    AND3 un13_nsum_adj_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[6] ));
    MX2 \LED_1[3]  (.A(LED_12_3), .B(LED_15_3), .S(choose_0_0), .Y(
        N_100));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I147_Y (.A(N535), .B(N531), 
        .Y(N596));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I121_Y (.A(N505), .B(N509), 
        .Y(N570));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I272_Y_0 (.A(
        ADD_32x32_fast_I272_un1_Y_0), .B(N638), .C(N637), .Y(
        ADD_32x32_fast_I272_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I173_Y (.A(N562), .B(N570), 
        .Y(N628));
    MX2 \sum_adj_RNO[9]  (.A(sum_9), .B(I_26_2), .S(sum_0_0), .Y(
        \nsum_adj_11[9] ));
    XA1 \off_div_RNO[22]  (.A(N767), .B(ADD_32x32_fast_I312_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[22] ));
    XOR2 \sum_adj_RNISADK[14]  (.A(\sum_adj[14]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[6] ));
    DFN1E1C0 \sum_adj[23]  (.D(\nsum_adj_11[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[23]_net_1 ));
    XOR2 \sum_adj_RNIO6DK[10]  (.A(\sum_adj[10]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[2] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I203_Y (.A(N594), .B(N601), 
        .C(N593), .Y(N659));
    NOR2 un13_nsum_adj_I_57 (.A(sum_18), .B(sum_19), .Y(
        \DWACT_FINC_E[14] ));
    XOR2 \sum_adj_RNIQ8DK[12]  (.A(\sum_adj[12]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[4] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I86_Y (.A(N389), .B(N393), .C(
        N392), .Y(N532));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I200_Y (.A(N597), .B(N590), 
        .C(N589), .Y(N655));
    MX2 \sum_adj_RNO[15]  (.A(sum_15), .B(I_43_2), .S(sum_2_0), .Y(
        \nsum_adj_11[15] ));
    NOR2A \LED_4[2]  (.A(LED_FB_2), .B(choose_0_0), .Y(N_52));
    XNOR2 un13_nsum_adj_I_53 (.A(sum_18), .B(N_7), .Y(I_53_2));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I315_Y_0 (.A(off_div[25]), 
        .B(sum_39), .Y(ADD_32x32_fast_I315_Y_0));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I84_Y (.A(N392), .B(
        off_div[4]), .C(\un1_sum_adj[4] ), .Y(N530));
    NOR3B un13_nsum_adj_I_45 (.A(\DWACT_FINC_E[10] ), .B(
        \DWACT_FINC_E[6] ), .C(sum_15), .Y(N_9));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I130_Y (.A(N518), .B(N515), 
        .C(N514), .Y(N579));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I118_Y (.A(N506), .B(N503), 
        .C(N502), .Y(N567));
    NOR3A \off_div_RNIJ6RC1[21]  (.A(next_off_div_2_sqmuxa_2), .B(
        off_div[21]), .C(off_div[23]), .Y(next_off_div_2_sqmuxa_6));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I273_un1_Y_0 (.A(N590), .B(
        N598), .C(\un1_sum_adj[0] ), .Y(ADD_32x32_fast_I273_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I69_Y (.A(N420), .B(N417), 
        .Y(N515));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I202_Y (.A(N592), .B(N599), 
        .C(N591), .Y(N657));
    NOR3C \off_div_RNITDOC1[17]  (.A(off_div[18]), .B(off_div[17]), .C(
        un5lto20_1), .Y(un5lto20_2));
    MX2 \sum_adj_RNO[16]  (.A(sum_16), .B(I_46_2), .S(sum_2_0), .Y(
        \nsum_adj_11[16] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I309_Y_0 (.A(off_div[19]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I309_Y_0));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I5_P0N (.A(sum_1_0), .B(
        \sum_adj[13]_net_1 ), .C(off_div[5]), .Y(N399));
    MX2 \off_div_RNO[3]  (.A(next_off_div_0_sqmuxa), .B(
        \un1_off_div_1[3] ), .S(\state_d_0[2] ), .Y(\next_off_div[3] ));
    AND3 un13_nsum_adj_I_69 (.A(\DWACT_FINC_E[29] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[33] ), .Y(N_2));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I76_Y (.A(N404), .B(N408), .C(
        N407), .Y(N522));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I4_G0N (.A(\un1_sum_adj[4] )
        , .B(off_div[4]), .Y(N395));
    NOR3A \off_div_RNIAC1D1[15]  (.A(un1_off_divlto31_8), .B(
        off_div[15]), .C(off_div[17]), .Y(un1_off_divlto31_15));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I1_P0N (.A(sum_1_0), .B(
        \sum_adj[9]_net_1 ), .C(off_div[1]), .Y(N387));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I13_G0N (.A(
        \un1_sum_adj[13] ), .B(off_div[13]), .Y(N422));
    DFN1E0C0 \off_div[15]  (.D(\next_off_div[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[15]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I150_Y (.A(I150_un1_Y), .B(
        N534), .Y(N599));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I144_Y (.A(N532), .B(N529), 
        .C(N528), .Y(N593));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I74_Y (.A(N407), .B(
        off_div[9]), .C(\un1_sum_adj[9] ), .Y(N520));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I50_Y (.A(off_div[20]), .B(
        off_div[21]), .C(sum_1_0), .Y(N496));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0_0 (.A(off_div[30]), 
        .B(off_div[29]), .C(sum_0_0), .Y(ADD_32x32_fast_I258_Y_0_0));
    DFN1E0C0 \off_div[13]  (.D(\next_off_div[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[13]));
    MX2 \sum_adj_RNO[20]  (.A(sum_20), .B(I_59_2), .S(sum_2_0), .Y(
        \nsum_adj_11[20] ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I293_Y_0 (.A(sum_2_0), .B(
        \sum_adj[11]_net_1 ), .C(off_div[3]), .Y(
        ADD_32x32_fast_I293_Y_0));
    AND2 un13_nsum_adj_I_44 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[9] ), .Y(\DWACT_FINC_E[10] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I272_un1_Y_0 (.A(N538), .B(
        N654), .Y(ADD_32x32_fast_I272_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I265_un1_Y (.A(
        ADD_32x32_fast_I265_un1_Y_0), .B(N802), .Y(I265_un1_Y));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I319_Y_0 (.A(off_div[29]), 
        .B(sum_39), .Y(ADD_32x32_fast_I319_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0_a3_0_1 (.A(N491), 
        .B(N487), .Y(ADD_32x32_fast_I258_Y_0_a3_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I265_Y_0 (.A(N557), .B(N565), 
        .Y(ADD_32x32_fast_I265_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I179_Y (.A(N568), .B(N576), 
        .Y(N634));
    AND3 un13_nsum_adj_I_39 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[8] ), .Y(N_11));
    XOR2 \sum_adj_RNI0FDK[18]  (.A(\sum_adj[18]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[10] ));
    XA1 \off_div_RNO[24]  (.A(N763), .B(ADD_32x32_fast_I314_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[24] ));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I309_Y (.A(I234_un1_Y), .B(
        ADD_32x32_fast_I270_Y_1), .C(ADD_32x32_fast_I309_Y_0), .Y(
        \un1_off_div_1[19] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0_a5_1 (.A(
        ADD_32x32_fast_I258_Y_0_a5_0), .B(N483), .Y(
        ADD_32x32_fast_I258_Y_0_a5_1));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I177_Y (.A(N566), .B(N574), 
        .Y(N632));
    OR2 \off_div_RNI1UVM[8]  (.A(off_div[8]), .B(off_div[9]), .Y(
        un5lto9));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I51_Y (.A(off_div[20]), .B(
        off_div[21]), .C(sum_1_0), .Y(N497));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I308_Y_0 (.A(off_div[18]), 
        .B(sum_39), .Y(ADD_32x32_fast_I308_Y_0));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I2_P0N (.A(sum_2_0), .B(
        \sum_adj[10]_net_1 ), .C(off_div[2]), .Y(N390));
    DFN1E0P0 \off_div[7]  (.D(\next_off_div[7] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2), .Q(off_div[7]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I196_Y (.A(I196_un1_Y), .B(
        N585), .Y(N651));
    NOR3 un13_nsum_adj_I_29 (.A(sum_7), .B(sum_6), .C(sum_8), .Y(
        \DWACT_FINC_E[5] ));
    XNOR2 un13_nsum_adj_I_65 (.A(sum_22), .B(N_3), .Y(I_65_2));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I268_Y (.A(I230_un1_Y), .B(
        N629), .C(I268_un1_Y), .Y(N769));
    DFN1E0C0 \off_div[9]  (.D(\next_off_div[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[9]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I37_Y (.A(off_div[27]), .B(
        off_div[28]), .C(sum_0_0), .Y(N483));
    DFN1E0C0 \off_div[11]  (.D(\next_off_div[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[11]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I145_Y (.A(N533), .B(N529), 
        .Y(N594));
    DFN1E1C0 \sum_adj[18]  (.D(\nsum_adj_11[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[18]_net_1 ));
    MX2 un1_off_div_1_0_0_ADD_32x32_fast_I92_Y (.A(sum_2_0), .B(
        off_div[0]), .S(\sum_adj[8]_net_1 ), .Y(N538));
    XA1 \off_div_RNO[13]  (.A(N787), .B(ADD_32x32_fast_I303_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[13] ));
    NOR2 \off_div_RNI0QDM[25]  (.A(off_div[27]), .B(off_div[25]), .Y(
        un1_off_divlto31_2));
    MX2 \sum_adj_RNO[21]  (.A(sum_21), .B(I_62_2), .S(sum_2_0), .Y(
        \nsum_adj_11[21] ));
    MX2 \LED_7[5]  (.A(N_47), .B(N_71), .S(choose[0]), .Y(LED_c_5));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I318_Y_0 (.A(off_div[28]), 
        .B(sum_39), .Y(ADD_32x32_fast_I318_Y_0));
    XNOR2 un13_nsum_adj_I_35 (.A(sum_12), .B(N_13), .Y(I_35_2));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I191_Y (.A(N588), .B(N580), 
        .Y(N646));
    MX2 \sum_adj_RNO[22]  (.A(sum_22), .B(I_65_2), .S(sum_2_0), .Y(
        \nsum_adj_11[22] ));
    MX2 \off_div_RNO[15]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[15] ), .S(\state_d[2] ), .Y(\next_off_div[15] ));
    NOR2 \off_div_RNILCBM[10]  (.A(off_div[10]), .B(off_div[13]), .Y(
        un1_off_divlto31_10));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I14_P0N (.A(sum_0_0), .B(
        \sum_adj[22]_net_1 ), .C(off_div[14]), .Y(N426));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0_a3_0_0 (.A(N560), 
        .B(N568), .Y(ADD_32x32_fast_I258_Y_0_a3_0_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I122_Y (.A(N510), .B(N507), 
        .C(N506), .Y(N571));
    NOR2 \off_div_RNIRKDM[22]  (.A(off_div[22]), .B(off_div[25]), .Y(
        next_off_div_2_sqmuxa_2));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I89_Y (.A(N387), .B(N390), 
        .Y(N535));
    AND3 un13_nsum_adj_I_64 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[16] ), .Y(N_3));
    OA1 \off_div_RNIM14U3[10]  (.A(un5lto9), .B(un5lt9), .C(
        off_div[10]), .Y(un5lt14));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I265_Y (.A(I224_un1_Y), .B(
        ADD_32x32_fast_I265_Y_0), .C(I265_un1_Y), .Y(N763));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I181_Y (.A(N578), .B(N570), 
        .Y(N636));
    NOR2A un13_nsum_adj_I_25 (.A(\DWACT_FINC_E[4] ), .B(sum_8), .Y(
        N_16));
    DFN1E1C0 \sum_adj[9]  (.D(\nsum_adj_11[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[9]_net_1 ));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I60_Y (.A(N428), .B(sum_1_0), 
        .C(off_div[16]), .Y(N506));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I307_Y (.A(I238_un1_Y), .B(
        ADD_32x32_fast_I272_Y_0), .C(ADD_32x32_fast_I307_Y_0), .Y(
        \un1_off_div_1[17] ));
    AND3 un13_nsum_adj_I_51 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[28] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I174_Y (.A(N571), .B(N564), 
        .C(N563), .Y(N629));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I140_Y (.A(N528), .B(N525), 
        .C(N524), .Y(N589));
    DFN1E1C0 \sum_adj[11]  (.D(\nsum_adj_11[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[11]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y_1 (.A(N620), .B(N635), 
        .C(ADD_32x32_fast_I263_Y_0), .Y(ADD_32x32_fast_I263_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I246_Y (.A(N650), .B(N599), 
        .C(N649), .Y(N793));
    XA1 \off_div_RNO[27]  (.A(N_6), .B(ADD_32x32_fast_I317_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[27] ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I291_Y_0 (.A(sum_0_0), .B(
        \sum_adj[9]_net_1 ), .C(off_div[1]), .Y(
        ADD_32x32_fast_I291_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I249_un1_Y (.A(N590), .B(
        N598), .C(\un1_sum_adj[0] ), .Y(I249_un1_Y));
    AND3 un13_nsum_adj_I_48 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[11] ), .Y(N_8));
    DFN1E0C0 \off_div[25]  (.D(\next_off_div[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[25]));
    XA1 \off_div_RNO[1]  (.A(N538), .B(ADD_32x32_fast_I291_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[1] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I61_Y (.A(N432), .B(N429), 
        .Y(N507));
    NOR2B un13_nsum_adj_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_13));
    DFN1E1C0 \sum_adj[22]  (.D(\nsum_adj_11[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[22]_net_1 ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I79_Y (.A(off_div[6]), .B(
        \un1_sum_adj[6] ), .C(N405), .Y(N525));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I150_un1_Y (.A(N535), .B(
        N538), .Y(I150_un1_Y));
    DFN1E0C0 \off_div[23]  (.D(\next_off_div[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[23]));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I304_Y_0 (.A(sum_1_0), .B(
        \sum_adj[22]_net_1 ), .C(off_div[14]), .Y(
        ADD_32x32_fast_I304_Y_0));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I298_Y_0 (.A(off_div[8]), .B(
        \un1_sum_adj[8] ), .Y(ADD_32x32_fast_I298_Y_0));
    XA1 \off_div_RNO[9]  (.A(N799), .B(ADD_32x32_fast_I299_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[9] ));
    NOR3A \off_div_RNIPCKO1[12]  (.A(un1_off_divlto31_0), .B(
        off_div[12]), .C(un5lto9), .Y(un1_off_divlto31_17));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y_1 (.A(N622), .B(N637), 
        .C(ADD_32x32_fast_I264_Y_0), .Y(ADD_32x32_fast_I264_Y_1));
    GND GND_i (.Y(GND));
    AND3 un13_nsum_adj_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E[4] ));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0_o5_0 (.A(N490), .B(
        N486), .Y(ADD_32x32_fast_I258_Y_0_o5_0));
    DFN1E1C0 \sum_adj[14]  (.D(\nsum_adj_11[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[14]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I138_Y (.A(N526), .B(N523), 
        .C(N522), .Y(N587));
    XOR2 \sum_adj_RNIFAHP[8]  (.A(\sum_adj[8]_net_1 ), .B(sum_39), .Y(
        \un1_sum_adj[0] ));
    OR2B \off_div_RNI4FF21[5]  (.A(un5lto4), .B(off_div[5]), .Y(
        un1_off_divlt31));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y (.A(
        ADD_32x32_fast_I259_un1_Y_0), .B(N784), .C(
        ADD_32x32_fast_I259_Y_3), .Y(N751));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I43_Y (.A(off_div[25]), .B(
        off_div[24]), .C(sum_0_0), .Y(N489));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I123_Y (.A(N507), .B(N511), 
        .Y(N572));
    XOR2 \sum_adj_RNIVDDK[17]  (.A(\sum_adj[17]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[9] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I175_Y (.A(N564), .B(N572), 
        .Y(N630));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I106_Y (.A(N494), .B(N490), 
        .Y(N555));
    MX2 \sum_adj_RNO[10]  (.A(sum_10), .B(I_28_2), .S(sum_2_0), .Y(
        \nsum_adj_11[10] ));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I11_G0N (.A(sum_0_0), .B(
        \sum_adj[19]_net_1 ), .C(off_div[11]), .Y(N416));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I314_Y_0 (.A(off_div[24]), 
        .B(sum_39), .Y(ADD_32x32_fast_I314_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I271_un1_Y_0 (.A(N586), .B(
        N594), .C(N601), .Y(ADD_32x32_fast_I271_un1_Y_0));
    DFN1E0C0 \off_div[21]  (.D(\next_off_div[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[21]));
    XA1 \off_div_RNO[11]  (.A(N793), .B(ADD_32x32_fast_I301_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[11] ));
    MX2 \LED_1[5]  (.A(LED_12_5), .B(LED_15_5), .S(choose_0_0), .Y(
        N_102));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I42_Y (.A(off_div[24]), .B(
        off_div[25]), .C(sum_0_0), .Y(N488));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y (.A(
        ADD_32x32_fast_I263_un1_Y_0), .B(N796), .C(
        ADD_32x32_fast_I263_Y_1), .Y(N759));
    OR2 \off_div_RNIHAT6A[31]  (.A(un1_off_div), .B(off_div[31]), .Y(
        next_off_div37));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I248_Y (.A(N654), .B(N538), 
        .C(N653), .Y(N799));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I301_Y_0 (.A(sum_2_0), .B(
        \sum_adj[19]_net_1 ), .C(off_div[11]), .Y(
        ADD_32x32_fast_I301_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y (.A(
        ADD_32x32_fast_I260_un1_Y_0), .B(N787), .C(
        ADD_32x32_fast_I260_Y_2), .Y(N753));
    AND3 un13_nsum_adj_I_68 (.A(\DWACT_FINC_E[34] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[29] ));
    NOR2A \LED_4[0]  (.A(LED_FB_0), .B(choose_0_0), .Y(N_50));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I306_Y_0 (.A(off_div[16]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I306_Y_0));
    NOR2 \off_div_RNISMEM[30]  (.A(off_div[27]), .B(off_div[30]), .Y(
        next_off_div_2_sqmuxa_4));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I80_Y (.A(N398), .B(
        off_div[6]), .C(\un1_sum_adj[6] ), .Y(N526));
    NOR3A \off_div_RNI3NRC1[26]  (.A(un1_off_divlto31_2), .B(
        off_div[26]), .C(off_div[29]), .Y(un1_off_divlto31_12));
    DFN1E1C0 \sum_adj[13]  (.D(\nsum_adj_11[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[13]_net_1 ));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I265_un1_Y_0 (.A(N582), .B(
        N574), .C(N624), .Y(ADD_32x32_fast_I265_un1_Y_0));
    NOR3C \state_RNIAO6TA[0]  (.A(state[1]), .B(state[0]), .C(
        next_off_div37), .Y(next_off_div_0_sqmuxa));
    DFN1E0C0 \off_div[5]  (.D(\next_off_div[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[5]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I7_G0N (.A(\un1_sum_adj[7] )
        , .B(off_div[7]), .Y(N404));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I57_Y (.A(off_div[17]), .B(
        off_div[18]), .C(sum_1_0), .Y(N503));
    XOR2 \state_RNO[1]  (.A(state[0]), .B(state[1]), .Y(N_311_i));
    OR2 \off_div_RNIPGBM[14]  (.A(off_div[14]), .B(off_div[13]), .Y(
        un5lto14_1));
    NOR3 un13_nsum_adj_I_18 (.A(sum_4), .B(sum_3), .C(sum_5), .Y(
        \DWACT_FINC_E[2] ));
    OR2 \off_div_RNINJVM[3]  (.A(off_div[4]), .B(off_div[3]), .Y(
        un5lto4));
    NOR2A \LED_5[0]  (.A(LED_33_0), .B(choose_0_0), .Y(N_58));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I308_Y (.A(I236_un1_Y), .B(
        ADD_32x32_fast_I271_Y_0), .C(ADD_32x32_fast_I308_Y_0), .Y(
        \un1_off_div_1[18] ));
    MX2 \sum_adj_RNO[11]  (.A(sum_11), .B(I_32_2), .S(sum_2_0), .Y(
        \nsum_adj_11[11] ));
    NOR3A \off_div_RNIH4RC1[23]  (.A(un1_off_divlto31_4), .B(
        off_div[23]), .C(off_div[24]), .Y(un1_off_divlto31_13));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I321_Y_0 (.A(off_div[31]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I321_Y_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I116_Y (.A(N504), .B(N500), 
        .Y(N565));
    NOR2 un13_nsum_adj_I_38 (.A(sum_12), .B(sum_13), .Y(
        \DWACT_FINC_E[8] ));
    AO1C \state_RNIQEBRL[1]  (.A(un5lt31), .B(next_off_div_2_sqmuxa_10)
        , .C(state[1]), .Y(un1_state_2));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I311_Y_0 (.A(off_div[21]), 
        .B(sum_39), .Y(ADD_32x32_fast_I311_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I269_Y_0 (.A(N647), .B(N632), 
        .C(N631), .Y(ADD_32x32_fast_I269_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I242_un1_Y_0 (.A(N584), .B(
        N576), .Y(ADD_32x32_fast_I242_un1_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I81_Y (.A(off_div[6]), .B(
        \un1_sum_adj[6] ), .C(N399), .Y(N527));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I245_Y (.A(N648), .B(N663), 
        .C(N647), .Y(N790));
    MX2 \sum_adj_RNO[12]  (.A(sum_12), .B(I_35_2), .S(sum_2_0), .Y(
        \nsum_adj_11[12] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I316_Y_0 (.A(off_div[26]), 
        .B(sum_39), .Y(ADD_32x32_fast_I316_Y_0));
    XNOR2 un13_nsum_adj_I_46 (.A(sum_16), .B(N_9), .Y(I_46_2));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I70_Y (.A(N413), .B(N417), .C(
        N416), .Y(N516));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I192_Y (.A(N589), .B(N582), 
        .C(N581), .Y(N647));
    XNOR2 un13_nsum_adj_I_28 (.A(sum_10), .B(N_15), .Y(I_28_2));
    NOR3A \off_div_RNITDOC1[19]  (.A(un1_off_divlto31_6), .B(
        off_div[19]), .C(off_div[21]), .Y(un1_off_divlto31_14));
    DFN1E0C0 \off_div[30]  (.D(\next_off_div[30] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[30]));
    NOR2 \off_div_RNI0OBM[16]  (.A(off_div[18]), .B(off_div[16]), .Y(
        un1_off_divlto31_6));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I129_Y (.A(N513), .B(N517), 
        .Y(N578));
    OA1 \off_div_RNIR5F21[1]  (.A(off_div[0]), .B(off_div[1]), .C(
        off_div[2]), .Y(un5lt4));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I182_Y (.A(N579), .B(N572), 
        .C(N571), .Y(N637));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I127_Y (.A(N511), .B(N515), 
        .Y(N576));
    VCC VCC_i (.Y(VCC));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I249_Y (.A(I249_un1_Y), .B(
        N655), .Y(N802));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I0_G0N (.A(off_div[0]), .B(
        sum_39), .Y(N383));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I196_un1_Y (.A(N593), .B(
        N586), .Y(I196_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I45_Y (.A(off_div[23]), .B(
        off_div[24]), .C(sum_1_0), .Y(N491));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I270_Y_1 (.A(
        ADD_32x32_fast_I270_un1_Y_0), .B(N599), .C(
        ADD_32x32_fast_I270_Y_0), .Y(ADD_32x32_fast_I270_Y_1));
    AND3 un13_nsum_adj_I_52 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[12] ), .Y(N_7));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I111_Y (.A(N495), .B(N499), 
        .Y(N560));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I71_Y (.A(N414), .B(N417), 
        .Y(N517));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I9_G0N (.A(\un1_sum_adj[9] )
        , .B(off_div[9]), .Y(N410));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I228_un1_Y (.A(N643), .B(
        N628), .Y(I228_un1_Y));
    MX2 \LED_3[0]  (.A(N_97), .B(N_34), .S(choose[1]), .Y(N_42));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I307_Y_0 (.A(off_div[17]), 
        .B(sum_39), .Y(ADD_32x32_fast_I307_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I2_G0N (.A(\un1_sum_adj[2] )
        , .B(off_div[2]), .Y(N389));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I148_Y (.A(N536), .B(N533), 
        .C(N532), .Y(N597));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I48_Y (.A(off_div[21]), .B(
        off_div[22]), .C(sum_1_0), .Y(N494));
    NOR2B \off_div_RNILGLR9[12]  (.A(un1_off_divlto31_22), .B(
        un1_off_divlto31_21), .Y(un1_off_div));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I260_un1_Y_0 (.A(N614), .B(
        N630), .Y(ADD_32x32_fast_I260_un1_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I268_un1_Y (.A(N630), .B(
        N646), .C(N661), .Y(I268_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_3 (.A(N612), .B(N627), 
        .C(ADD_32x32_fast_I259_Y_2), .Y(ADD_32x32_fast_I259_Y_3));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0_o5 (.A(
        ADD_32x32_fast_I258_Y_0_a3_0), .B(N_5), .C(
        ADD_32x32_fast_I258_Y_0_o5_0), .Y(N_6));
    NOR3C \off_div_RNI88A95[15]  (.A(un1_off_divlto31_15), .B(
        un1_off_divlto31_14), .C(un1_off_divlto31_20), .Y(
        un1_off_divlto31_22));
    NOR2A \LED_2[0]  (.A(LED_5_0), .B(choose[2]), .Y(N_34));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I67_Y (.A(off_div[13]), .B(
        \un1_sum_adj[13] ), .C(N420), .Y(N513));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0_o3_0 (.A(N494), .B(
        N498), .Y(ADD_32x32_fast_I258_Y_0_o3_0));
    XNOR2 un13_nsum_adj_I_70 (.A(sum_23), .B(N_2), .Y(I_70_2));
    NOR3A un13_nsum_adj_I_66 (.A(\DWACT_FINC_E[15] ), .B(sum_21), .C(
        sum_22), .Y(\DWACT_FINC_E[33] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I193_Y (.A(N582), .B(N590), 
        .Y(N648));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I5_G0N (.A(sum_1_0), .B(
        \sum_adj[13]_net_1 ), .C(off_div[5]), .Y(N398));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I317_Y_0 (.A(off_div[27]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I317_Y_0));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y_1 (.A(N482), .B(N486), 
        .C(N555), .Y(ADD_32x32_fast_I260_Y_1));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0_1 (.A(
        ADD_32x32_fast_I258_Y_0_0), .B(N482), .Y(
        ADD_32x32_fast_I258_Y_0_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I243_Y (.A(N644), .B(N659), 
        .C(N643), .Y(N784));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I296_Y_0 (.A(off_div[6]), .B(
        \un1_sum_adj[6] ), .Y(ADD_32x32_fast_I296_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I183_Y (.A(N572), .B(N580), 
        .Y(N638));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I157_Y_1 (.A(
        ADD_32x32_fast_I157_Y_0), .B(N485), .Y(ADD_32x32_fast_I157_Y_1)
        );
    MX2 \sum_adj_RNO[8]  (.A(sum_8), .B(I_23_8), .S(sum_0_0), .Y(
        \nsum_adj_11[8] ));
    XA1 \off_div_RNO[6]  (.A(N659), .B(ADD_32x32_fast_I296_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[6] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I124_Y (.A(N512), .B(N509), 
        .C(N508), .Y(N573));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I157_Y_0 (.A(off_div[29]), .B(
        off_div[28]), .C(sum_0_0), .Y(ADD_32x32_fast_I157_Y_0));
    NOR3C \off_div_RNID8BI4[12]  (.A(un1_off_divlto31_13), .B(
        un1_off_divlto31_12), .C(un1_off_divlto31_17), .Y(
        un1_off_divlto31_21));
    NOR3B un13_nsum_adj_I_36 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .C(sum_12), .Y(N_12));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I242_Y (.A(
        ADD_32x32_fast_I242_un1_Y_0), .B(N657), .C(
        ADD_32x32_fast_I242_Y_0), .Y(N781));
    NOR3C \off_div_RNIALF21[5]  (.A(off_div[6]), .B(off_div[7]), .C(
        off_div[5]), .Y(un5lto7_1));
    DFN1E0C0 \off_div[1]  (.D(\next_off_div[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[1]));
    NOR2 un13_nsum_adj_I_47 (.A(sum_15), .B(sum_16), .Y(
        \DWACT_FINC_E[11] ));
    XA1 \off_div_RNO[8]  (.A(N802), .B(ADD_32x32_fast_I298_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[8] ));
    XNOR2 un13_nsum_adj_I_26 (.A(sum_9), .B(N_16), .Y(I_26_2));
    XOR2 \sum_adj_RNISBEK[23]  (.A(\sum_adj[23]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[15] ));
    XNOR2 un13_nsum_adj_I_43 (.A(sum_15), .B(N_10), .Y(I_43_2));
    NOR2B \off_div_RNISKCM[19]  (.A(off_div[20]), .B(off_div[19]), .Y(
        un5lto20_1));
    MX2 \off_div_RNO[19]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[19] ), .S(\state_d[2] ), .Y(\next_off_div[19] ));
    DFN1E0C0 \off_div[10]  (.D(\next_off_div[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[10]));
    MX2 \off_div_RNO[10]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[10] ), .S(\state_d[2] ), .Y(\next_off_div[10] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I125_Y (.A(N513), .B(N509), 
        .Y(N574));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y_0 (.A(N553), .B(N561), 
        .Y(ADD_32x32_fast_I263_Y_0));
    NOR3C \off_div_RNIUAAR3[21]  (.A(next_off_div_2_sqmuxa_6), .B(
        next_off_div_2_sqmuxa_5), .C(next_off_div_2_sqmuxa_7), .Y(
        next_off_div_2_sqmuxa_9));
    DFN1E1C0 \sum_adj[12]  (.D(\nsum_adj_11[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[12]_net_1 ));
    NOR3 un13_nsum_adj_I_50 (.A(sum_15), .B(sum_17), .C(sum_16), .Y(
        \DWACT_FINC_E[12] ));
    MX2 \sum_adj_RNO[17]  (.A(sum_17), .B(I_49_2), .S(sum_2_0), .Y(
        \nsum_adj_11[17] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0_o3_1 (.A(N560), .B(
        N567), .C(ADD_32x32_fast_I258_Y_0_o3_0), .Y(
        ADD_32x32_fast_I258_Y_0_o3_1));
    NOR2A \LED_5[2]  (.A(LED_33_2), .B(choose_0_0), .Y(N_60));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I297_Y (.A(\un1_sum_adj[7] ), 
        .B(off_div[7]), .C(N657), .Y(\un1_off_div_1[7] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I269_un1_Y (.A(
        ADD_32x32_fast_I269_un1_Y_0), .B(N663), .Y(I269_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I136_Y (.A(N524), .B(N521), 
        .C(N520), .Y(N585));
    XA1 \off_div_RNO[16]  (.A(N779), .B(ADD_32x32_fast_I306_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[16] ));
    MX2 \off_div_RNO[0]  (.A(next_off_div_0_sqmuxa), .B(
        \un1_off_div_1[0] ), .S(\state_d_0[2] ), .Y(\next_off_div[0] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I199_Y (.A(N596), .B(N588), 
        .Y(N654));
    XA1 \off_div_RNO[23]  (.A(N_5), .B(ADD_32x32_fast_I313_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[23] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I264_un1_Y_0 (.A(N622), .B(
        N638), .Y(ADD_32x32_fast_I264_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I87_Y (.A(N390), .B(N393), 
        .Y(N533));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I189_Y (.A(N578), .B(N586), 
        .Y(N644));
    MX2 \off_div_RNO[18]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[18] ), .S(\state_d[2] ), .Y(\next_off_div[18] ));
    MX2 \LED_6[0]  (.A(N_50), .B(N_58), .S(choose[1]), .Y(N_66));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I38_Y (.A(off_div[27]), .B(
        off_div[26]), .C(sum_0_0), .Y(N484));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I273_Y (.A(I273_un1_Y), .B(
        N639), .C(I240_un1_Y), .Y(N779));
    NOR3 un13_nsum_adj_I_67 (.A(sum_0_d0), .B(sum_2_d0), .C(sum_1_d0), 
        .Y(\DWACT_FINC_E[34] ));
    XA1 \off_div_RNO[25]  (.A(N761), .B(ADD_32x32_fast_I315_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[25] ));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I112_Y (.A(N496), .B(N500), 
        .Y(N561));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I14_G0N (.A(sum_0_0), .B(
        \sum_adj[22]_net_1 ), .C(off_div[14]), .Y(N425));
    XOR2 \sum_adj_RNIUCDK[16]  (.A(\sum_adj[16]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[8] ));
    DFN1E0C0 \off_div[12]  (.D(\next_off_div[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[12]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I271_Y_0 (.A(
        ADD_32x32_fast_I271_un1_Y_0), .B(N636), .C(N635), .Y(
        ADD_32x32_fast_I271_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0_o3 (.A(
        ADD_32x32_fast_I258_Y_0_a3_0_0), .B(N781), .C(
        ADD_32x32_fast_I258_Y_0_o3_1), .Y(N_5));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I161_Y (.A(N485), .B(N489), 
        .C(N558), .Y(N616));
    DFN1E0C0 \off_div[0]  (.D(\next_off_div[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[0]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I234_un1_Y (.A(N634), .B(
        N649), .Y(I234_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I131_Y (.A(N515), .B(N519), 
        .Y(N580));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I120_Y (.A(N508), .B(N505), 
        .C(N504), .Y(N569));
    NOR2A un13_nsum_adj_I_63 (.A(\DWACT_FINC_E[15] ), .B(sum_21), .Y(
        \DWACT_FINC_E[16] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I46_Y (.A(off_div[22]), .B(
        off_div[23]), .C(sum_1_0), .Y(N492));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I300_Y_0 (.A(off_div[10]), 
        .B(\un1_sum_adj[10] ), .Y(ADD_32x32_fast_I300_Y_0));
    NOR2 \off_div_RNI8ILM[11]  (.A(off_div[6]), .B(off_div[11]), .Y(
        un1_off_divlto31_9));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I77_Y (.A(N405), .B(N408), 
        .Y(N523));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I44_Y (.A(off_div[23]), .B(
        off_div[24]), .C(sum_0_0), .Y(N490));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y_2 (.A(N614), .B(N629), 
        .C(ADD_32x32_fast_I260_Y_1), .Y(ADD_32x32_fast_I260_Y_2));
    DFN1E1C0 \sum_adj[20]  (.D(\nsum_adj_11[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[20]_net_1 ));
    NOR2A \LED_2[3]  (.A(LED_5_3), .B(choose[2]), .Y(N_37));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I53_Y (.A(off_div[20]), .B(
        off_div[19]), .C(sum_1_0), .Y(N499));
    MX2 \off_div_RNO[5]  (.A(next_off_div_0_sqmuxa), .B(
        \un1_off_div_1[5] ), .S(\state_d_0[2] ), .Y(\next_off_div[5] ));
    XNOR2 un13_nsum_adj_I_37 (.A(sum_13), .B(N_12), .Y(I_37_2));
    XA1 \off_div_RNO[2]  (.A(N601), .B(ADD_32x32_fast_I292_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[2] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I6_G0N (.A(\un1_sum_adj[6] )
        , .B(off_div[6]), .Y(N401));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I247_un1_Y (.A(N586), .B(
        N594), .C(N601), .Y(I247_un1_Y));
    NOR3B \state_RNIAO6TA_0[0]  (.A(state[1]), .B(state[0]), .C(
        next_off_div37), .Y(next_off_div_1_sqmuxa));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I151_Y (.A(N537), .B(
        \un1_sum_adj[0] ), .C(N536), .Y(N601));
    DFN1E0C0 \off_div[6]  (.D(\next_off_div[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[6]));
    NOR3 un13_nsum_adj_I_33 (.A(sum_10), .B(sum_9), .C(sum_11), .Y(
        \DWACT_FINC_E[7] ));
    DFN1E1C0 \sum_adj[17]  (.D(\nsum_adj_11[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[17]_net_1 ));
    NOR2 \off_div_RNICMLM[14]  (.A(off_div[14]), .B(off_div[7]), .Y(
        un1_off_divlto31_8));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I320_Y_0 (.A(off_div[30]), 
        .B(sum_39), .Y(ADD_32x32_fast_I320_Y_0));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I305_Y (.A(\un1_sum_adj[15] )
        , .B(off_div[15]), .C(N781), .Y(\un1_off_div_1[15] ));
    NOR3A un13_nsum_adj_I_27 (.A(\DWACT_FINC_E[4] ), .B(sum_8), .C(
        sum_9), .Y(N_15));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I310_Y_0 (.A(off_div[20]), 
        .B(sum_39), .Y(ADD_32x32_fast_I310_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I270_Y_0 (.A(N575), .B(N568), 
        .C(N567), .Y(ADD_32x32_fast_I270_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I230_un1_Y (.A(N645), .B(
        N630), .Y(I230_un1_Y));
    NOR2A \LED_4[5]  (.A(LED_FB_5), .B(choose_0_0), .Y(N_55));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I52_Y (.A(off_div[20]), .B(
        off_div[19]), .C(sum_1_0), .Y(N498));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I204_Y (.A(I204_un1_Y), .B(
        N595), .Y(N661));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I263_un1_Y_0 (.A(N620), .B(
        N636), .Y(ADD_32x32_fast_I263_un1_Y_0));
    MX2 \LED_3[2]  (.A(N_99), .B(N_36), .S(choose[1]), .Y(N_44));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I194_Y (.A(N591), .B(N584), 
        .C(N583), .Y(N649));
    XNOR2 un13_nsum_adj_I_23 (.A(sum_8), .B(N_17), .Y(I_23_8));
    NOR2A \LED_2[5]  (.A(LED_5_5), .B(choose[2]), .Y(N_39));
    XNOR2 un13_nsum_adj_I_59 (.A(sum_20), .B(N_5_0), .Y(I_59_2));
    DFN1E0C0 \off_div[20]  (.D(\next_off_div[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[20]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I113_Y (.A(N501), .B(N497), 
        .Y(N562));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I184_Y (.A(N581), .B(N574), 
        .C(N573), .Y(N639));
    NOR3 un13_nsum_adj_I_41 (.A(sum_13), .B(sum_12), .C(sum_14), .Y(
        \DWACT_FINC_E[9] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_0 (.A(off_div[28]), .B(
        off_div[29]), .C(sum_2_0), .Y(ADD_32x32_fast_I259_Y_0));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I294_Y_0 (.A(off_div[4]), .B(
        \un1_sum_adj[4] ), .Y(ADD_32x32_fast_I294_Y_0));
    MX2 \LED_6[5]  (.A(N_55), .B(N_63), .S(choose[1]), .Y(N_71));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I236_un1_Y (.A(N651), .B(
        N636), .Y(I236_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I10_G0N (.A(
        \un1_sum_adj[10] ), .B(off_div[10]), .Y(N413));
    XA1 \off_div_RNO[21]  (.A(N769), .B(ADD_32x32_fast_I311_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[21] ));
    DFN1E0C0 \off_div[18]  (.D(\next_off_div[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[18]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I109_Y (.A(N497), .B(N493), 
        .Y(N558));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I146_Y (.A(N534), .B(N531), 
        .C(N530), .Y(N595));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I107_Y (.A(N495), .B(N491), 
        .Y(N556));
    OA1 \off_div_RNISEUR2[1]  (.A(un5lto4), .B(un5lt4), .C(un5lto7_1), 
        .Y(un5lt9));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I195_Y (.A(N592), .B(N584), 
        .Y(N650));
    NOR2 \off_div_RNIMFDM[20]  (.A(off_div[22]), .B(off_div[20]), .Y(
        un1_off_divlto31_4));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I63_Y (.A(N429), .B(N426), 
        .Y(N509));
    NOR3B un13_nsum_adj_I_55 (.A(\DWACT_FINC_E[13] ), .B(
        \DWACT_FINC_E[28] ), .C(sum_18), .Y(N_6_0));
    DFN1E0C0 \off_div[22]  (.D(\next_off_div[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[22]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I90_Y (.A(N383), .B(N387), .C(
        N386), .Y(N536));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I55_Y (.A(off_div[18]), .B(
        off_div[19]), .C(sum_1_0), .Y(N501));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I49_Y (.A(off_div[22]), .B(
        off_div[21]), .C(sum_1_0), .Y(N495));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_2 (.A(N484), .B(
        ADD_32x32_fast_I259_Y_0), .C(N553), .Y(ADD_32x32_fast_I259_Y_2)
        );
    XA1 \off_div_RNO[12]  (.A(N790), .B(ADD_32x32_fast_I302_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[12] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I62_Y (.A(N425), .B(N429), .C(
        N428), .Y(N508));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y (.A(
        ADD_32x32_fast_I261_un1_Y_0), .B(N790), .C(
        ADD_32x32_fast_I261_Y_2), .Y(N755));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I141_Y (.A(N529), .B(N525), 
        .Y(N590));
    AND3 un13_nsum_adj_I_61 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[15] ), .Y(N_4));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I36_Y (.A(off_div[28]), .B(
        off_div[27]), .C(sum_0_0), .Y(N482));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I7_P0N (.A(\un1_sum_adj[7] ), 
        .B(off_div[7]), .Y(N405));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I58_Y (.A(off_div[17]), .B(
        off_div[16]), .C(sum_1_0), .Y(N504));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I292_Y_0 (.A(off_div[2]), .B(
        \un1_sum_adj[2] ), .Y(ADD_32x32_fast_I292_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I91_Y (.A(sum_1_0), .B(
        off_div[0]), .C(N387), .Y(N537));
    DFN1E0C0 \off_div[17]  (.D(\next_off_div[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[17]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I119_Y (.A(N503), .B(N507), 
        .Y(N568));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I190_Y (.A(N587), .B(N580), 
        .C(N579), .Y(N645));
    AND3 un13_nsum_adj_I_54 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[9] ), .C(\DWACT_FINC_E[12] ), .Y(
        \DWACT_FINC_E[13] ));
    MX2 \sum_adj_RNO[23]  (.A(sum_23), .B(I_70_2), .S(sum_2_0), .Y(
        \nsum_adj_11[23] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I117_Y (.A(N501), .B(N505), 
        .Y(N566));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I132_Y (.A(N520), .B(N517), 
        .C(N516), .Y(N581));
    OA1 \off_div_RNI2P0M5[15]  (.A(un5lt14), .B(un5lto14_2), .C(
        off_div[15]), .Y(un5lt16));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I180_Y (.A(N577), .B(N570), 
        .C(N569), .Y(N635));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I128_Y (.A(N516), .B(N513), 
        .C(N512), .Y(N577));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I104_Y (.A(N492), .B(N488), 
        .Y(N553));
    NOR3A un13_nsum_adj_I_31 (.A(\DWACT_FINC_E[6] ), .B(sum_9), .C(
        sum_10), .Y(N_14));
    XOR2 \sum_adj_RNIQ9EK[21]  (.A(\sum_adj[21]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[13] ));
    OA1 \off_div_RNIU1VD7[16]  (.A(off_div[16]), .B(un5lt16), .C(
        un5lto20_2), .Y(un5lt31));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I240_un1_Y (.A(N582), .B(
        N574), .C(N655), .Y(I240_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I15_G0N (.A(
        \un1_sum_adj[15] ), .B(off_div[15]), .Y(N428));
    NOR2 \off_div_RNITNEM[30]  (.A(off_div[30]), .B(off_div[28]), .Y(
        un1_off_divlto31_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I273_un1_Y (.A(N582), .B(
        N574), .C(ADD_32x32_fast_I273_un1_Y_0), .Y(I273_un1_Y));
    NOR2 un13_nsum_adj_I_21 (.A(sum_6), .B(sum_7), .Y(
        \DWACT_FINC_E[3] ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I295_Y_0 (.A(sum_0_0), .B(
        \sum_adj[13]_net_1 ), .C(off_div[5]), .Y(
        ADD_32x32_fast_I295_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I176_Y (.A(N573), .B(N566), 
        .C(N565), .Y(N631));
    DFN1E0C0 \off_div[28]  (.D(\next_off_div[28] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[28]));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I83_Y (.A(off_div[4]), .B(
        \un1_sum_adj[4] ), .C(N399), .Y(N529));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I65_Y (.A(off_div[13]), .B(
        \un1_sum_adj[13] ), .C(N426), .Y(N511));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I12_P0N (.A(sum_1_0), .B(
        \sum_adj[20]_net_1 ), .C(off_div[12]), .Y(N420));
    DFN1C0 \state[1]  (.D(N_311_i), .CLK(clk_c), .CLR(n_rst_c), .Q(
        state[1]));
    MX2 \LED_3[3]  (.A(N_100), .B(N_37), .S(choose[1]), .Y(N_45));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I15_P0N (.A(\un1_sum_adj[15] )
        , .B(off_div[15]), .Y(N429));
    XA1 \off_div_RNO[31]  (.A(N749), .B(ADD_32x32_fast_I321_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[31] ));
    XA1 \off_div_RNO[14]  (.A(N784), .B(ADD_32x32_fast_I304_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[14] ));
    MX2 \LED_7[0]  (.A(N_42), .B(N_66), .S(choose[0]), .Y(LED_c_0));
    AND3 un13_nsum_adj_I_42 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[9] ), .Y(N_10));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I133_Y (.A(N517), .B(N521), 
        .Y(N582));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I68_Y (.A(N416), .B(N420), .C(
        N419), .Y(N514));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I114_Y (.A(N502), .B(N498), 
        .Y(N563));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I261_un1_Y_0 (.A(N616), .B(
        N632), .Y(ADD_32x32_fast_I261_un1_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I82_Y (.A(N395), .B(N399), .C(
        N398), .Y(N528));
    MX2 \sum_adj_RNO[14]  (.A(sum_14), .B(I_40_2), .S(sum_2_0), .Y(
        \nsum_adj_11[14] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I40_Y (.A(off_div[25]), .B(
        off_div[26]), .C(sum_0_0), .Y(N486));
    DFN1E1C0 \sum_adj[8]  (.D(\nsum_adj_11[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[8]_net_1 ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I204_un1_Y (.A(N596), .B(
        N538), .Y(I204_un1_Y));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I12_G0N (.A(sum_1_0), .B(
        \sum_adj[20]_net_1 ), .C(off_div[12]), .Y(N419));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I11_P0N (.A(sum_0_0), .B(
        \sum_adj[19]_net_1 ), .C(off_div[11]), .Y(N417));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I73_Y (.A(off_div[9]), .B(
        \un1_sum_adj[9] ), .C(N414), .Y(N519));
    MX2 \LED_1[2]  (.A(LED_12_2), .B(LED_15_2), .S(choose_0_0), .Y(
        N_99));
    AO1C \state_RNIQEBRL_0[1]  (.A(un5lt31), .B(
        next_off_div_2_sqmuxa_10), .C(state[1]), .Y(un1_state_2_0));
    MX2 \LED_1[0]  (.A(LED_12_0), .B(LED_15_0), .S(choose_0_0), .Y(
        N_97));
    AND3 un13_nsum_adj_I_58 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[14] ), .Y(N_5_0));
    OA1B \state_RNO[0]  (.A(state[1]), .B(pwm_enable), .C(state[0]), 
        .Y(\state_ns[0] ));
    DFN1E0C0 \off_div[2]  (.D(\next_off_div[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[2]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I39_Y (.A(off_div[26]), .B(
        off_div[27]), .C(sum_0_0), .Y(N485));
    DFN1E0C0 \off_div[27]  (.D(\next_off_div[27] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[27]));
    MX2 \sum_adj_RNO[18]  (.A(sum_18), .B(I_53_2), .S(sum_2_0), .Y(
        \nsum_adj_11[18] ));
    DFN1E1C0 \sum_adj[15]  (.D(\nsum_adj_11[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[15]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I41_Y (.A(off_div[26]), .B(
        off_div[25]), .C(sum_0_0), .Y(N487));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y (.A(
        ADD_32x32_fast_I264_un1_Y_0), .B(N799), .C(
        ADD_32x32_fast_I264_Y_1), .Y(N761));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I72_Y (.A(N410), .B(N414), .C(
        N413), .Y(N518));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I295_Y (.A(
        ADD_32x32_fast_I295_Y_0), .B(N661), .Y(\un1_off_div_1[5] ));
    XA1 \off_div_RNO[29]  (.A(N753), .B(ADD_32x32_fast_I319_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[29] ));
    DFN1E0C0 \off_div[14]  (.D(\next_off_div[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[14]));
    DFN1E1C0 \sum_adj[10]  (.D(\nsum_adj_11[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[10]_net_1 ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I302_Y_0 (.A(sum_0_0), .B(
        \sum_adj[20]_net_1 ), .C(off_div[12]), .Y(
        ADD_32x32_fast_I302_Y_0));
    MX2 \off_div_RNO[20]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[20] ), .S(\state_d[2] ), .Y(\next_off_div[20] ));
    OR3 \off_div_RNIETMC1[11]  (.A(off_div[11]), .B(off_div[12]), .C(
        un5lto14_1), .Y(un5lto14_2));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I300_Y (.A(
        ADD_32x32_fast_I300_Y_0), .B(N796), .Y(\un1_off_div_1[10] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I115_Y (.A(N499), .B(N503), 
        .Y(N564));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I142_Y (.A(N530), .B(N527), 
        .C(N526), .Y(N591));
    XNOR2 un13_nsum_adj_I_62 (.A(sum_21), .B(N_4), .Y(I_62_2));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I56_Y (.A(off_div[17]), .B(
        off_div[18]), .C(sum_1_0), .Y(N502));
    XA1 \off_div_RNO[26]  (.A(N759), .B(ADD_32x32_fast_I316_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[26] ));
    MX2 \sum_adj_RNO[13]  (.A(sum_13), .B(I_37_2), .S(sum_2_0), .Y(
        \nsum_adj_11[13] ));
    DFN1E1C0 \sum_adj[19]  (.D(\nsum_adj_11[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[19]_net_1 ));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I267_un1_Y (.A(N628), .B(
        N644), .C(N659), .Y(I267_un1_Y));
    MX2 \off_div_RNO[17]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[17] ), .S(\state_d[2] ), .Y(\next_off_div[17] ));
    NOR2A \state_RNIPD9M_1[0]  (.A(state[0]), .B(state[1]), .Y(
        state_176_d));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I54_Y (.A(off_div[18]), .B(
        off_div[19]), .C(sum_1_0), .Y(N500));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I267_Y (.A(I228_un1_Y), .B(
        N627), .C(I267_un1_Y), .Y(N767));
    DFN1E0P0 \off_div[4]  (.D(\next_off_div[4] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2), .Q(off_div[4]));
    NOR2A \LED_5[5]  (.A(LED_33_5), .B(choose[2]), .Y(N_63));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I303_Y_0 (.A(off_div[13]), 
        .B(\un1_sum_adj[13] ), .Y(ADD_32x32_fast_I303_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I169_Y (.A(N566), .B(N558), 
        .Y(N624));
    DFN1E0C0 \off_div[19]  (.D(\next_off_div[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[19]));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I85_Y (.A(off_div[4]), .B(
        \un1_sum_adj[4] ), .C(N393), .Y(N531));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I312_Y_0 (.A(off_div[22]), 
        .B(sum_39), .Y(ADD_32x32_fast_I312_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I270_un1_Y_0 (.A(N650), .B(
        N634), .Y(ADD_32x32_fast_I270_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I139_Y (.A(N527), .B(N523), 
        .Y(N588));
    XA1 \off_div_RNO[28]  (.A(N755), .B(ADD_32x32_fast_I318_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[28] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I167_Y (.A(N556), .B(N564), 
        .Y(N622));
    DFN1E0C0 \off_div[16]  (.D(\next_off_div[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[16]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I8_P0N (.A(\un1_sum_adj[8] ), 
        .B(off_div[8]), .Y(N408));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I198_Y (.A(N595), .B(N588), 
        .C(N587), .Y(N653));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I137_Y (.A(N525), .B(N521), 
        .Y(N586));
    DFN1E0P0 \off_div[8]  (.D(\next_off_div[8] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2), .Q(off_div[8]));
    XNOR2 un13_nsum_adj_I_32 (.A(sum_11), .B(N_14), .Y(I_32_2));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I188_Y (.A(N585), .B(N578), 
        .C(N577), .Y(N643));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I16_P0N (.A(off_div[16]), .B(
        sum_39), .Y(N432));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I88_Y (.A(N386), .B(N390), .C(
        N389), .Y(N534));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0 (.A(
        ADD_32x32_fast_I258_Y_0_a5_1), .B(N_6), .C(
        ADD_32x32_fast_I258_Y_0_1), .Y(N749));
    AND3 un13_nsum_adj_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_17));
    XOR2 \sum_adj_RNITBDK[15]  (.A(\sum_adj[15]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[7] ));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I310_Y (.A(I269_un1_Y), .B(
        ADD_32x32_fast_I269_Y_0), .C(ADD_32x32_fast_I310_Y_0), .Y(
        \un1_off_div_1[20] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y_2 (.A(N616), .B(N631), 
        .C(ADD_32x32_fast_I261_Y_1), .Y(ADD_32x32_fast_I261_Y_2));
    NOR3C \off_div_RNI1EGF2[10]  (.A(un1_off_divlto31_10), .B(
        un1_off_divlto31_9), .C(un1_off_divlt31), .Y(
        un1_off_divlto31_20));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I159_Y (.A(N483), .B(N487), 
        .C(N556), .Y(N614));
    XNOR2 un13_nsum_adj_I_40 (.A(sum_14), .B(N_11), .Y(I_40_2));
    NOR3A \off_div_RNIUISC1[26]  (.A(next_off_div_2_sqmuxa_4), .B(
        off_div[28]), .C(off_div[26]), .Y(next_off_div_2_sqmuxa_7));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I242_Y_0 (.A(N583), .B(N576), 
        .C(N575), .Y(ADD_32x32_fast_I242_Y_0));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I313_Y_0 (.A(off_div[23]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I313_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I157_Y (.A(N489), .B(N493), 
        .C(ADD_32x32_fast_I157_Y_1), .Y(N612));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I75_Y (.A(off_div[9]), .B(
        \un1_sum_adj[9] ), .C(N408), .Y(N521));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I293_Y (.A(
        ADD_32x32_fast_I293_Y_0), .B(N599), .Y(\un1_off_div_1[3] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I143_Y (.A(N531), .B(N527), 
        .Y(N592));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I259_un1_Y_0 (.A(N612), .B(
        N628), .Y(ADD_32x32_fast_I259_un1_Y_0));
    DFN1E0C0 \off_div[3]  (.D(\next_off_div[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2), .Q(off_div[3]));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I290_Y (.A(sum_0_0), .B(
        off_div[0]), .C(\un1_sum_adj[0] ), .Y(\un1_off_div_1[0] ));
    XNOR2 un13_nsum_adj_I_56 (.A(sum_19), .B(N_6_0), .Y(I_56_2));
    MX2 \off_div_RNO[7]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[7] ), .S(\state_d_0[2] ), .Y(\next_off_div[7] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I78_Y (.A(N401), .B(N405), .C(
        N404), .Y(N524));
    DFN1E1C0 \sum_adj[21]  (.D(\nsum_adj_11[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[21]_net_1 ));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I66_Y (.A(N419), .B(
        off_div[13]), .C(\un1_sum_adj[13] ), .Y(N512));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I8_G0N (.A(\un1_sum_adj[8] )
        , .B(off_div[8]), .Y(N407));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I224_un1_Y (.A(N624), .B(
        N639), .Y(I224_un1_Y));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I299_Y_0 (.A(off_div[9]), .B(
        \un1_sum_adj[9] ), .Y(ADD_32x32_fast_I299_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I269_un1_Y_0 (.A(N648), .B(
        N632), .Y(ADD_32x32_fast_I269_un1_Y_0));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I1_G0N (.A(sum_1_0), .B(
        \sum_adj[9]_net_1 ), .C(off_div[1]), .Y(N386));
    XA1 \off_div_RNO[4]  (.A(N663), .B(ADD_32x32_fast_I294_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[4] ));
    DFN1E0C0 \off_div[24]  (.D(\next_off_div[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[24]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0_a5_0 (.A(off_div[29])
        , .B(off_div[30]), .C(sum_0_0), .Y(
        ADD_32x32_fast_I258_Y_0_a5_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I64_Y (.A(N422), .B(N426), .C(
        N425), .Y(N510));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I205_Y (.A(N598), .B(
        \un1_sum_adj[0] ), .C(N597), .Y(N663));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I172_Y (.A(N569), .B(N562), 
        .C(N561), .Y(N627));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I3_G0N (.A(sum_0_0), .B(
        \sum_adj[11]_net_1 ), .C(off_div[3]), .Y(N392));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I134_Y (.A(N522), .B(N519), 
        .C(N518), .Y(N583));
    DFN1E1C0 \sum_adj[16]  (.D(\nsum_adj_11[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[16]_net_1 ));
    MX2 \LED_3[5]  (.A(N_102), .B(N_39), .S(choose[1]), .Y(N_47));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I244_Y (.A(N646), .B(N661), 
        .C(N645), .Y(N787));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I238_un1_Y (.A(N653), .B(
        N638), .Y(I238_un1_Y));
    MX2 \LED_7[2]  (.A(N_44), .B(N_68), .S(choose[0]), .Y(LED_c_2));
    MX2 \sum_adj_RNO[19]  (.A(sum_19), .B(I_56_2), .S(sum_2_0), .Y(
        \nsum_adj_11[19] ));
    NOR2A \state_RNIPD9M_0[0]  (.A(state[1]), .B(state[0]), .Y(
        \state_d[2] ));
    NOR2A \off_div_RNIFL72E[31]  (.A(next_off_div_2_sqmuxa_9), .B(
        next_off_div37), .Y(next_off_div_2_sqmuxa_10));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y_1 (.A(N484), .B(N488), 
        .C(N557), .Y(ADD_32x32_fast_I261_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I126_Y (.A(N514), .B(N511), 
        .C(N510), .Y(N575));
    NOR3 un13_nsum_adj_I_60 (.A(sum_19), .B(sum_18), .C(sum_20), .Y(
        \DWACT_FINC_E[15] ));
    XA1 \off_div_RNO[30]  (.A(N751), .B(ADD_32x32_fast_I320_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[30] ));
    
endmodule


module integral_calc_13s_4_2(
       avg_old,
       avg_new,
       LED_5,
       average,
       LED_5_i_0,
       calc_avg,
       avg_done,
       n_rst_c,
       clk_c
    );
input  [11:0] avg_old;
input  [11:0] avg_new;
output [7:0] LED_5;
output [6:2] average;
output LED_5_i_0;
input  calc_avg;
output avg_done;
input  n_rst_c;
input  clk_c;

    wire \state_1[0]_net_1 , \state_1_RNIQNJE[0]_net_1 , 
        \state_0[0]_net_1 , avg_done_0, \state[1]_net_1 , 
        ADD_26x26_fast_I253_Y_0, \integ[23]_net_1 , 
        ADD_26x26_fast_I254_Y_0, \integ[24]_net_1 , \state[0]_net_1 , 
        ADD_26x26_fast_I255_Y_0, \integ[25]_net_1 , 
        ADD_26x26_fast_I206_Y_2, N506, N521, ADD_26x26_fast_I206_Y_1, 
        N402, N398, N459, ADD_26x26_fast_I252_Y_0, \integ[22]_net_1 , 
        ADD_26x26_fast_I204_Y_3, N517, N502, ADD_26x26_fast_I204_Y_2, 
        ADD_26x26_fast_I204_Y_0, N455, ADD_26x26_fast_I205_Y_3, N504, 
        N519, ADD_26x26_fast_I205_Y_2, ADD_26x26_fast_I205_Y_1, N457, 
        ADD_26x26_fast_I205_Y_0, N400, ADD_26x26_fast_I250_Y_0, 
        \integ[20]_net_1 , ADD_26x26_fast_I251_Y_0, \integ[21]_net_1 , 
        ADD_26x26_fast_I249_Y_0, \integ[19]_net_1 , 
        ADD_26x26_fast_I207_Y_2, N508, N523, ADD_26x26_fast_I207_Y_1, 
        N404, N461, ADD_26x26_fast_I246_Y_0, \integ[16]_net_1 , 
        ADD_26x26_fast_I248_Y_0, \integ[18]_net_1 , 
        ADD_26x26_fast_I247_Y_0, \integ[17]_net_1 , 
        ADD_26x26_fast_I241_Y_0, \un1_next_int[11] , 
        ADD_26x26_fast_I209_Y_1, ADD_26x26_fast_I209_un1_Y_0, N543, 
        ADD_26x26_fast_I209_Y_0, N465, N458, ADD_26x26_fast_I208_Y_1, 
        ADD_26x26_fast_I208_un1_Y_0, N541, ADD_26x26_fast_I208_Y_0, 
        N456, N463, ADD_26x26_fast_I238_Y_0, \un1_next_int[8] , 
        ADD_26x26_fast_I239_Y_0, \un18_next_int_m[9] , \inf_abs0_m[9] , 
        ADD_26x26_fast_I210_Y_1, ADD_26x26_fast_I210_un1_Y_0, N491, 
        ADD_26x26_fast_I210_Y_0, N467, N460, 
        ADD_26x26_fast_I204_un1_Y_0, N518, ADD_26x26_fast_I205_un1_Y_0, 
        N520, ADD_26x26_fast_I240_Y_0, \un1_next_int[10] , 
        ADD_26x26_fast_I213_Y_0, ADD_26x26_fast_I213_un1_Y_0, 
        ADD_26x26_fast_I211_Y_1, ADD_26x26_fast_I211_un1_Y_0, N532, 
        ADD_26x26_fast_I211_Y_0, N469, N462, ADD_26x26_fast_I212_Y_0, 
        ADD_26x26_fast_I212_un1_Y_0, ADD_26x26_fast_I234_Y_0, 
        \state_RNIFCE11[0]_net_1 , ADD_26x26_fast_I235_Y_0, 
        \un1_next_int[5] , N510, N526, N512, N528, N476, N484, N514, 
        N480, N488, N442, N482, N490, \state_RNI74E11[0]_net_1 , N470, 
        N493, ADD_26x26_fast_I232_Y_0, \state_RNIB8E11[0]_net_1 , 
        ADD_26x26_fast_I231_Y_0, \inf_abs0_m[1] , \un18_next_int_m[1] , 
        \integ[1]_net_1 , ADD_26x26_fast_I125_Y_0, 
        ADD_26x26_fast_I127_Y_0, ADD_26x26_fast_I230_Y_0, 
        \integ[0]_net_1 , ADD_26x26_fast_I230_Y_1, \un1_integ[11] , 
        N529, I192_un1_Y, N401, N405, I205_un1_Y, N535, I195_un1_Y, 
        I207_un1_Y, N524, N539, N403, N399, I206_un1_Y, N522, N537, 
        \un1_integ[22] , \un1_integ[23] , \un1_integ[3] , 
        \un1_next_int[3] , \un1_integ[24] , \un1_integ[16] , 
        I186_un1_Y, \un1_integ[17] , I184_un1_Y, \un1_integ[15] , 
        \integ[15]_net_1 , N637, I204_un1_Y, N533, I194_un1_Y, 
        \un1_integ[4] , \un1_integ[8] , \un1_integ[20] , I178_un1_Y, 
        \un1_integ[25] , \un1_integ[10] , N531, I193_un1_Y, 
        \un1_integ[5] , \un1_integ[6] , \un1_next_int[6] , 
        \un1_integ[19] , I180_un1_Y, \un1_integ[18] , I182_un1_Y, 
        \un1_integ[14] , N640, \un1_integ[2] , \un1_integ[12] , N646, 
        \un1_integ[7] , \state_RNILIE11[0]_net_1 , \un1_integ[13] , 
        N643, \un1_integ[21] , I176_un1_Y, \un1_integ[9] , 
        \un1_integ[1] , N527, N423, N348, N345, N525, N422, N344, N347, 
        N413, N415, N357, N477, N428, N425, N424, N478, N429, N409, 
        N412, N408, N486, N485, \inf_abs0_m[10] , 
        \un18_next_int_m[10] , N436, N433, N432, N437, I110_un1_Y, 
        N481, N416, N466, N417, N421, N354, N353, N420, N474, N473, 
        N414, N411, N410, N407, N406, N341, I152_un1_Y, N475, N483, 
        N468, N342, I150_un1_Y, I163_un1_Y, N489, \inf_abs0_m[11] , 
        \un18_next_int_m[11] , N418, N350, N351, N419, N487, N479, 
        N430, N427, N426, N439, N324, N321, N464, N472, N471, N441, 
        N318, N338, I74_un1_Y, N317, N438, I148_un1_Y, N320, N323, 
        N440, \inf_abs0_m[3] , \un18_next_int_m[3] , \inf_abs0_m[4] , 
        \un18_next_int_m[4] , \inf_abs0_m[7] , \un18_next_int_m[7] , 
        \inf_abs0_m[2] , \un18_next_int_m[2] , \inf_abs0_m[5] , 
        \un18_next_int_m[5] , \inf_abs0_m[6] , \un18_next_int_m[6] , 
        N336, N332, I121_un1_Y, I64_un1_Y, N329, N333, N330, N327, 
        N326, N434, N335, N435, N431, \state_RNO_5[1] , I162_un1_Y, 
        I112_un1_Y, \inf_abs0_m[0] , \un18_next_int_m[0] , 
        \inf_abs0_m[8] , \un18_next_int_m[8] , GND, VCC;
    
    AO1 un1_integ_0_0_ADD_26x26_fast_I56_Y (.A(N341), .B(N345), .C(
        N344), .Y(N424));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I148_un1_Y (.A(N479), .B(N472), 
        .Y(I148_un1_Y));
    DFN1C0 \state[0]  (.D(\state_1_RNIQNJE[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state[0]_net_1 ));
    DFN1E0C0 \integ[13]  (.D(\un1_integ[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_5[6]));
    NOR2B \state_RNINVAG[0]  (.A(avg_new[6]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[6] ));
    DFN1E0C0 \integ[24]  (.D(\un1_integ[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[24]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I112_un1_Y (.A(N434), .B(N431), 
        .Y(I112_un1_Y));
    OA1 un1_integ_0_0_ADD_26x26_fast_I61_Y (.A(
        \state_RNILIE11[0]_net_1 ), .B(LED_5[0]), .C(N336), .Y(N429));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I248_Y_0 (.A(\integ[18]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I248_Y_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I41_Y (.A(\integ[16]_net_1 ), .B(
        \integ[17]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N409));
    NOR2B \state_RNIO0BG[0]  (.A(avg_new[7]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[7] ));
    NOR2B \state_RNIKSAG[0]  (.A(avg_new[3]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[3] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I204_un1_Y (.A(N533), .B(
        I194_un1_Y), .C(ADD_26x26_fast_I204_un1_Y_0), .Y(I204_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I86_Y (.A(N408), .B(N404), .Y(
        N457));
    AO1 un1_integ_0_0_ADD_26x26_fast_I98_Y (.A(N420), .B(N417), .C(
        N416), .Y(N469));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I176_un1_Y (.A(N525), .B(N510), 
        .Y(I176_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I205_un1_Y_0 (.A(N504), .B(N520)
        , .Y(ADD_26x26_fast_I205_un1_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I150_un1_Y (.A(N481), .B(N474), 
        .Y(I150_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I51_Y (.A(N354), .B(N351), .Y(
        N419));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y (.A(
        ADD_26x26_fast_I230_Y_0), .B(\state_RNI74E11[0]_net_1 ), .Y(
        ADD_26x26_fast_I230_Y_1));
    AX1D un1_integ_0_0_ADD_26x26_fast_I253_Y (.A(I206_un1_Y), .B(
        ADD_26x26_fast_I206_Y_2), .C(ADD_26x26_fast_I253_Y_0), .Y(
        \un1_integ[23] ));
    DFN1E0C0 \integ[21]  (.D(\un1_integ[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[21]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I146_Y (.A(N477), .B(N470), .C(
        N469), .Y(N523));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I210_un1_Y_0 (.A(N476), .B(N484)
        , .C(N514), .Y(ADD_26x26_fast_I210_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I142_Y (.A(N473), .B(N466), .C(
        N465), .Y(N519));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I231_Y (.A(
        ADD_26x26_fast_I231_Y_0), .B(N442), .Y(\un1_integ[1] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I155_Y (.A(N486), .B(N478), .Y(
        N532));
    DFN1E0C0 \integ[15]  (.D(\un1_integ[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[15]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I103_Y (.A(N421), .B(N425), .Y(
        N474));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I125_Y (.A(N399), .B(
        ADD_26x26_fast_I125_Y_0), .C(N456), .Y(N502));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_1 (.A(
        ADD_26x26_fast_I209_un1_Y_0), .B(N543), .C(
        ADD_26x26_fast_I209_Y_0), .Y(ADD_26x26_fast_I209_Y_1));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I97_Y (.A(N415), .B(N419), .Y(
        N468));
    NOR2B \state_RNIQ2BG[0]  (.A(avg_new[9]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[9] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I94_Y (.A(N416), .B(N413), .C(
        N412), .Y(N465));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I151_Y (.A(N482), .B(N474), .Y(
        N528));
    OR2 un1_integ_0_0_ADD_26x26_fast_I74_Y (.A(I74_un1_Y), .B(N317), 
        .Y(N442));
    AX1D un1_integ_0_0_ADD_26x26_fast_I238_Y (.A(N535), .B(I195_un1_Y), 
        .C(ADD_26x26_fast_I238_Y_0), .Y(\un1_integ[8] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I121_Y (.A(I121_un1_Y), .B(N440), 
        .Y(N493));
    AO1 un1_integ_0_0_ADD_26x26_fast_I190_Y (.A(N526), .B(N541), .C(
        N525), .Y(N643));
    OR2 un1_integ_0_0_ADD_26x26_fast_I5_P0N (.A(average[5]), .B(
        \un1_next_int[5] ), .Y(N333));
    NOR2B \state_RNIP1BG[0]  (.A(avg_new[8]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[8] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I246_Y (.A(I186_un1_Y), .B(
        ADD_26x26_fast_I213_Y_0), .C(ADD_26x26_fast_I246_Y_0), .Y(
        \un1_integ[16] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I252_Y_0 (.A(\integ[22]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I252_Y_0));
    DFN1C0 \state_1[0]  (.D(\state_1_RNIQNJE[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_1[0]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I39_Y (.A(\integ[17]_net_1 ), .B(
        \integ[18]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N407));
    OA1B un1_integ_0_0_ADD_26x26_fast_I32_Y (.A(\integ[21]_net_1 ), .B(
        \integ[20]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N400));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I194_un1_Y (.A(N480), .B(N488), 
        .C(N442), .Y(I194_un1_Y));
    AO1B un1_integ_0_0_ADD_26x26_fast_I125_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\integ[24]_net_1 ), .C(\state_1[0]_net_1 ), .Y(
        ADD_26x26_fast_I125_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I100_Y (.A(N422), .B(N419), .C(
        N418), .Y(N471));
    OR2 un1_integ_0_0_ADD_26x26_fast_I12_P0N (.A(LED_5[5]), .B(
        \state[1]_net_1 ), .Y(N354));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I10_G0N (.A(\un1_next_int[10] ), 
        .B(LED_5[3]), .Y(N347));
    DFN1E0C0 \integ[12]  (.D(\un1_integ[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_5[5]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I109_Y (.A(N427), .B(N431), .Y(
        N480));
    OR2 \state_RNIFCE11[0]  (.A(\inf_abs0_m[4] ), .B(
        \un18_next_int_m[4] ), .Y(\state_RNIFCE11[0]_net_1 ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I205_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\integ[22]_net_1 ), .C(\state_1[0]_net_1 ), .Y(
        ADD_26x26_fast_I205_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I115_Y (.A(N437), .B(N433), .Y(
        N486));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I12_G0N (.A(LED_5[5]), .B(
        \state[1]_net_1 ), .Y(N353));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_0 (.A(N456), .B(N463), .C(
        N455), .Y(ADD_26x26_fast_I208_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I111_Y (.A(N433), .B(N429), .Y(
        N482));
    OR2 un1_integ_0_0_ADD_26x26_fast_I2_P0N (.A(average[2]), .B(
        \state_RNIB8E11[0]_net_1 ), .Y(N324));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I250_Y_0 (.A(\integ[20]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I250_Y_0));
    DFN1E0C0 \integ[10]  (.D(\un1_integ[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_5[3]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I180_un1_Y (.A(N514), .B(N529), 
        .Y(I180_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I162_Y (.A(I162_un1_Y), .B(N487), 
        .Y(N541));
    NOR2A \state_RNIVJ3H[1]  (.A(\state[1]_net_1 ), .B(avg_old[9]), .Y(
        \un18_next_int_m[9] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I6_G0N (.A(average[6]), .B(
        \un1_next_int[6] ), .Y(N335));
    AX1D un1_integ_0_0_ADD_26x26_fast_I249_Y (.A(I180_un1_Y), .B(
        ADD_26x26_fast_I210_Y_1), .C(ADD_26x26_fast_I249_Y_0), .Y(
        \un1_integ[19] ));
    GND GND_i (.Y(GND));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I246_Y_0 (.A(\integ[16]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I246_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I6_P0N (.A(average[6]), .B(
        \un1_next_int[6] ), .Y(N336));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I212_un1_Y_0 (.A(N480), .B(N488)
        , .C(N442), .Y(ADD_26x26_fast_I212_un1_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I1_G0N (.A(\inf_abs0_m[1] ), .B(
        \un18_next_int_m[1] ), .C(\integ[1]_net_1 ), .Y(N320));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I107_Y (.A(N429), .B(N425), .Y(
        N478));
    OA1B un1_integ_0_0_ADD_26x26_fast_I38_Y (.A(\integ[17]_net_1 ), .B(
        \integ[18]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N406));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I209_un1_Y_0 (.A(N512), .B(N528)
        , .Y(ADD_26x26_fast_I209_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_3 (.A(N504), .B(N519), .C(
        ADD_26x26_fast_I205_Y_2), .Y(ADD_26x26_fast_I205_Y_3));
    AX1D un1_integ_0_0_ADD_26x26_fast_I255_Y (.A(I204_un1_Y), .B(
        ADD_26x26_fast_I204_Y_3), .C(ADD_26x26_fast_I255_Y_0), .Y(
        \un1_integ[25] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I204_Y_0 (.A(\integ[24]_net_1 ), 
        .B(\integ[23]_net_1 ), .C(\state_0[0]_net_1 ), .Y(
        ADD_26x26_fast_I204_Y_0));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I243_Y (.A(\state_0[0]_net_1 ), 
        .B(LED_5[6]), .C(N643), .Y(\un1_integ[13] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I231_Y_0 (.A(\inf_abs0_m[1] ), 
        .B(\un18_next_int_m[1] ), .C(\integ[1]_net_1 ), .Y(
        ADD_26x26_fast_I231_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I69_Y (.A(N327), .B(N324), .Y(
        N437));
    AO1 un1_integ_0_0_ADD_26x26_fast_I62_Y (.A(N332), .B(N336), .C(
        N335), .Y(N430));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I193_un1_Y (.A(N532), .B(N493), 
        .Y(I193_un1_Y));
    NOR2A \state_RNIUI3H[1]  (.A(\state[1]_net_1 ), .B(avg_old[8]), .Y(
        \un18_next_int_m[8] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I152_un1_Y (.A(N476), .B(N483), 
        .Y(I152_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I7_G0N (.A(LED_5[0]), .B(
        \state_RNILIE11[0]_net_1 ), .Y(N338));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I49_Y (.A(N354), .B(N357), .Y(
        N417));
    OA1B un1_integ_0_0_ADD_26x26_fast_I42_Y (.A(\integ[15]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_1[0]_net_1 ), .Y(N410));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I145_Y (.A(N468), .B(N476), .Y(
        N522));
    OR2 un1_integ_0_0_ADD_26x26_fast_I10_P0N (.A(\un1_next_int[10] ), 
        .B(LED_5[3]), .Y(N348));
    INV \integ_RNIFMD7[12]  (.A(LED_5[5]), .Y(LED_5_i_0));
    NOR2A \state_RNISG3H[1]  (.A(\state[1]_net_1 ), .B(avg_old[6]), .Y(
        \un18_next_int_m[6] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I1_P0N (.A(\inf_abs0_m[1] ), .B(
        \un18_next_int_m[1] ), .C(\integ[1]_net_1 ), .Y(N321));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I184_un1_Y (.A(N533), .B(N518), 
        .Y(I184_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I192_un1_Y (.A(N476), .B(N484), 
        .C(N491), .Y(I192_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I141_Y (.A(N464), .B(N472), .Y(
        N518));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I93_Y (.A(N411), .B(N415), .Y(
        N464));
    AO1B un1_integ_0_0_ADD_26x26_fast_I37_Y (.A(\integ[19]_net_1 ), .B(
        \integ[18]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N405));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I0_G0N (.A(\integ[0]_net_1 ), 
        .B(\state[1]_net_1 ), .Y(N317));
    OR2 \state_RNIPQHK[1]  (.A(\un18_next_int_m[10] ), .B(
        \inf_abs0_m[10] ), .Y(\un1_next_int[10] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I73_Y (.A(N318), .B(N321), .Y(
        N441));
    OA1 un1_integ_0_0_ADD_26x26_fast_I59_Y (.A(
        \state_RNILIE11[0]_net_1 ), .B(LED_5[0]), .C(N342), .Y(N427));
    AO1 un1_integ_0_0_ADD_26x26_fast_I52_Y (.A(N347), .B(N351), .C(
        N350), .Y(N420));
    NOR2A \state_RNO[1]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 ), 
        .Y(\state_RNO_5[1] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I34_Y (.A(\integ[20]_net_1 ), .B(
        \integ[19]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N402));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I236_Y (.A(\un1_next_int[6] ), 
        .B(average[6]), .C(N539), .Y(\un1_integ[6] ));
    NOR2B \state_RNIJRAG[0]  (.A(avg_new[2]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[2] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I205_Y_1 (.A(
        ADD_26x26_fast_I205_Y_0), .B(N400), .Y(ADD_26x26_fast_I205_Y_1)
        );
    OR2 un1_integ_0_0_ADD_26x26_fast_I150_Y (.A(I150_un1_Y), .B(N473), 
        .Y(N527));
    DFN1C0 \integ[0]  (.D(ADD_26x26_fast_I230_Y_1), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\integ[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I120_Y (.A(N439), .B(N442), .C(
        N438), .Y(N491));
    AO1 un1_integ_0_0_ADD_26x26_fast_I104_Y (.A(N426), .B(N423), .C(
        N422), .Y(N475));
    VCC VCC_i (.Y(VCC));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I129_Y (.A(N403), .B(N399), .C(
        N460), .Y(N506));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I113_Y (.A(N431), .B(N435), .Y(
        N484));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I241_Y_0 (.A(LED_5[4]), .B(
        \un1_next_int[11] ), .Y(ADD_26x26_fast_I241_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I89_Y (.A(N411), .B(N407), .Y(
        N460));
    AO1 un1_integ_0_0_ADD_26x26_fast_I68_Y (.A(N323), .B(N327), .C(
        N326), .Y(N436));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_0 (.A(N469), .B(N462), .C(
        N461), .Y(ADD_26x26_fast_I211_Y_0));
    DFN1E0C0 \integ[4]  (.D(\un1_integ[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[4]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I108_Y (.A(N430), .B(N427), .C(
        N426), .Y(N479));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I3_G0N (.A(average[3]), .B(
        \un1_next_int[3] ), .Y(N326));
    AO13 un1_integ_0_0_ADD_26x26_fast_I48_Y (.A(LED_5[6]), .B(N353), 
        .C(\state_1[0]_net_1 ), .Y(N416));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I195_un1_Y (.A(N482), .B(N490), 
        .C(\state_RNI74E11[0]_net_1 ), .Y(I195_un1_Y));
    DFN1E0C0 \integ[3]  (.D(\un1_integ[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[3]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I252_Y (.A(I207_un1_Y), .B(
        ADD_26x26_fast_I207_Y_2), .C(ADD_26x26_fast_I252_Y_0), .Y(
        \un1_integ[22] ));
    NOR2A \state_RNIOC3H[1]  (.A(\state[1]_net_1 ), .B(avg_old[2]), .Y(
        \un18_next_int_m[2] ));
    DFN1E0C0 \integ[6]  (.D(\un1_integ[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[6]));
    NOR2A \state_RNIMA3H[1]  (.A(\state[1]_net_1 ), .B(avg_old[0]), .Y(
        \un18_next_int_m[0] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_1 (.A(
        ADD_26x26_fast_I210_un1_Y_0), .B(N491), .C(
        ADD_26x26_fast_I210_Y_0), .Y(ADD_26x26_fast_I210_Y_1));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y (.A(N533), .B(I194_un1_Y), 
        .C(ADD_26x26_fast_I239_Y_0), .Y(\un1_integ[9] ));
    NOR2A \state_RNITH3H[1]  (.A(\state[1]_net_1 ), .B(avg_old[7]), .Y(
        \un18_next_int_m[7] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I58_Y (.A(N338), .B(N342), .C(
        N341), .Y(N426));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I67_Y (.A(N327), .B(N330), .Y(
        N435));
    OR2 \state_RNI74E11[0]  (.A(\un18_next_int_m[0] ), .B(
        \inf_abs0_m[0] ), .Y(\state_RNI74E11[0]_net_1 ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I253_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I253_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I64_Y (.A(I64_un1_Y), .B(N332), 
        .Y(N432));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I204_un1_Y_0 (.A(N502), .B(N518)
        , .Y(ADD_26x26_fast_I204_un1_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I127_Y (.A(N401), .B(
        ADD_26x26_fast_I127_Y_0), .C(N458), .Y(N504));
    OR2 un1_integ_0_0_ADD_26x26_fast_I110_Y (.A(I110_un1_Y), .B(N428), 
        .Y(N481));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I211_un1_Y_0 (.A(N470), .B(N462)
        , .C(N493), .Y(ADD_26x26_fast_I211_un1_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I90_Y (.A(N412), .B(N408), .Y(
        N461));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I233_Y (.A(\un1_next_int[3] ), 
        .B(average[3]), .C(N491), .Y(\un1_integ[3] ));
    OA1A un1_integ_0_0_ADD_26x26_fast_I47_Y (.A(\state_1[0]_net_1 ), 
        .B(LED_5[7]), .C(N357), .Y(N415));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I119_Y (.A(N441), .B(N437), .Y(
        N490));
    AO1 un1_integ_0_0_ADD_26x26_fast_I70_Y (.A(N320), .B(N324), .C(
        N323), .Y(N438));
    DFN1E0C0 \integ[5]  (.D(\un1_integ[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[5]));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I182_un1_Y (.A(N470), .B(N462), 
        .C(N531), .Y(I182_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I161_Y (.A(N486), .B(N493), .C(
        N485), .Y(N539));
    OA1B un1_integ_0_0_ADD_26x26_fast_I44_Y (.A(\integ[15]_net_1 ), .B(
        LED_5[7]), .C(\state_1[0]_net_1 ), .Y(N412));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I245_Y (.A(\state_0[0]_net_1 ), 
        .B(\integ[15]_net_1 ), .C(N637), .Y(\un1_integ[15] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I95_Y (.A(N417), .B(N413), .Y(
        N466));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y_0 (.A(
        \un18_next_int_m[9] ), .B(\inf_abs0_m[9] ), .C(LED_5[2]), .Y(
        ADD_26x26_fast_I239_Y_0));
    DFN1E0C0 \integ[2]  (.D(\un1_integ[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[2]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I135_Y (.A(N458), .B(N466), .Y(
        N512));
    OR2 un1_integ_0_0_ADD_26x26_fast_I88_Y (.A(N406), .B(N410), .Y(
        N459));
    AX1D un1_integ_0_0_ADD_26x26_fast_I247_Y (.A(I184_un1_Y), .B(
        ADD_26x26_fast_I212_Y_0), .C(ADD_26x26_fast_I247_Y_0), .Y(
        \un1_integ[17] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I143_Y (.A(N466), .B(N474), .Y(
        N520));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I57_Y (.A(N342), .B(N345), .Y(
        N425));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I186_un1_Y (.A(N535), .B(N520), 
        .Y(I186_un1_Y));
    DFN1E0C0 \integ[23]  (.D(\un1_integ[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[23]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I8_P0N (.A(\un1_next_int[8] ), .B(
        LED_5[1]), .Y(N342));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_2 (.A(N506), .B(N521), .C(
        ADD_26x26_fast_I206_Y_1), .Y(ADD_26x26_fast_I206_Y_2));
    AO1 un1_integ_0_0_ADD_26x26_fast_I54_Y (.A(N344), .B(N348), .C(
        N347), .Y(N422));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I131_Y (.A(N401), .B(N405), .C(
        N462), .Y(N508));
    OR2 \state_RNILIE11[0]  (.A(\inf_abs0_m[7] ), .B(
        \un18_next_int_m[7] ), .Y(\state_RNILIE11[0]_net_1 ));
    NOR2 \state_1_RNITM7C[0]  (.A(\state[1]_net_1 ), .B(
        \state_1[0]_net_1 ), .Y(avg_done));
    AX1D un1_integ_0_0_ADD_26x26_fast_I254_Y (.A(I205_un1_Y), .B(
        ADD_26x26_fast_I205_Y_3), .C(ADD_26x26_fast_I254_Y_0), .Y(
        \un1_integ[24] ));
    DFN1E0C0 \integ[19]  (.D(\un1_integ[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[19]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I117_Y (.A(N439), .B(N435), .Y(
        N488));
    OR2 \state_RNIDAE11[0]  (.A(\inf_abs0_m[3] ), .B(
        \un18_next_int_m[3] ), .Y(\un1_next_int[3] ));
    DFN1E0C0 \integ[17]  (.D(\un1_integ[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[17]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I33_Y (.A(\integ[20]_net_1 ), .B(
        \integ[21]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N401));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I255_Y_0 (.A(\integ[25]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I255_Y_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I127_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\integ[22]_net_1 ), .C(\state_0[0]_net_1 ), .Y(
        ADD_26x26_fast_I127_Y_0));
    DFN1E0C0 \integ[14]  (.D(\un1_integ[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_5[7]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I87_Y (.A(N405), .B(N409), .Y(
        N458));
    NOR2A \state_RNIPD3H[1]  (.A(\state[1]_net_1 ), .B(avg_old[3]), .Y(
        \un18_next_int_m[3] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y_0 (.A(average[2]), .B(
        \state_RNIB8E11[0]_net_1 ), .Y(ADD_26x26_fast_I232_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I84_Y (.A(N402), .B(N406), .Y(
        N455));
    AO1 un1_integ_0_0_ADD_26x26_fast_I154_Y (.A(N485), .B(N478), .C(
        N477), .Y(N531));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I11_G0N (.A(\un1_next_int[11] ), 
        .B(LED_5[4]), .Y(N350));
    AO1 un1_integ_0_0_ADD_26x26_fast_I140_Y (.A(N471), .B(N464), .C(
        N463), .Y(N517));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I149_Y (.A(N480), .B(N472), .Y(
        N526));
    AO1 un1_integ_0_0_ADD_26x26_fast_I158_Y (.A(N489), .B(N482), .C(
        N481), .Y(N535));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I249_Y_0 (.A(\integ[19]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I249_Y_0));
    DFN1E0C0 \integ[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[25]_net_1 ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I247_Y_0 (.A(\integ[17]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I247_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y_0 (.A(\integ[0]_net_1 ), 
        .B(\state[1]_net_1 ), .Y(ADD_26x26_fast_I230_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I64_un1_Y (.A(N329), .B(N333), 
        .Y(I64_un1_Y));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I242_Y (.A(\state[1]_net_1 ), .B(
        LED_5[5]), .C(N646), .Y(\un1_integ[12] ));
    DFN1E0C0 \integ[11]  (.D(\un1_integ[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_5[4]));
    DFN1E0C0 \integ[16]  (.D(\un1_integ[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[16]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_1 (.A(
        ADD_26x26_fast_I211_un1_Y_0), .B(N532), .C(
        ADD_26x26_fast_I211_Y_0), .Y(ADD_26x26_fast_I211_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I189_Y (.A(N524), .B(N539), .C(
        N523), .Y(N640));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I254_Y_0 (.A(\integ[24]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I254_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I163_Y (.A(I163_un1_Y), .B(N489), 
        .Y(N543));
    AO1 un1_integ_0_0_ADD_26x26_fast_I96_Y (.A(N418), .B(N415), .C(
        N414), .Y(N467));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I207_un1_Y (.A(N524), .B(N508), 
        .C(N539), .Y(I207_un1_Y));
    NOR2B \state_RNIIQAG[0]  (.A(avg_new[1]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[1] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I2_G0N (.A(average[2]), .B(
        \state_RNIB8E11[0]_net_1 ), .Y(N323));
    AO1 un1_integ_0_0_ADD_26x26_fast_I114_Y (.A(N436), .B(N433), .C(
        N432), .Y(N485));
    NOR2B \state_1_RNIJB8G[0]  (.A(avg_new[11]), .B(\state_1[0]_net_1 )
        , .Y(\inf_abs0_m[11] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I147_Y (.A(N470), .B(N478), .Y(
        N524));
    DFN1E0C0 \integ[9]  (.D(\un1_integ[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(LED_5[2]));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I235_Y (.A(
        ADD_26x26_fast_I235_Y_0), .B(N541), .Y(\un1_integ[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I212_Y_0 (.A(
        ADD_26x26_fast_I212_un1_Y_0), .B(N518), .C(N517), .Y(
        ADD_26x26_fast_I212_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I63_Y (.A(N333), .B(N336), .Y(
        N431));
    NOR2A \state_RNI8H94[1]  (.A(\state[1]_net_1 ), .B(avg_old[11]), 
        .Y(\un18_next_int_m[11] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I118_Y (.A(N440), .B(N437), .C(
        N436), .Y(N489));
    NOR2B \state_RNILTAG[0]  (.A(avg_new[4]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[4] ));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I237_Y (.A(
        \state_RNILIE11[0]_net_1 ), .B(LED_5[0]), .C(N537), .Y(
        \un1_integ[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I133_Y (.A(N456), .B(N464), .Y(
        N510));
    OA1B un1_integ_0_0_ADD_26x26_fast_I30_Y (.A(\integ[22]_net_1 ), .B(
        \integ[21]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N398));
    DFN1E0C0 \integ[22]  (.D(\un1_integ[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[22]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I43_Y (.A(\integ[15]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_1[0]_net_1 ), .Y(N411));
    DFN1E0C0 \integ[1]  (.D(\un1_integ[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(\integ[1]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I35_Y (.A(\integ[19]_net_1 ), .B(
        \integ[20]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N403));
    DFN1C0 \state_0[0]  (.D(\state_1_RNIQNJE[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_0[0]_net_1 ));
    OR2 \state_RNINKE11[0]  (.A(\un18_next_int_m[8] ), .B(
        \inf_abs0_m[8] ), .Y(\un1_next_int[8] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I53_Y (.A(N351), .B(N348), .Y(
        N421));
    AO1 un1_integ_0_0_ADD_26x26_fast_I160_Y (.A(N484), .B(N491), .C(
        N483), .Y(N537));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I91_Y (.A(N409), .B(N413), .Y(
        N462));
    AX1D un1_integ_0_0_ADD_26x26_fast_I250_Y (.A(I178_un1_Y), .B(
        ADD_26x26_fast_I209_Y_1), .C(ADD_26x26_fast_I250_Y_0), .Y(
        \un1_integ[20] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I240_Y_0 (.A(LED_5[3]), .B(
        \un1_next_int[10] ), .Y(ADD_26x26_fast_I240_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_0 (.A(N467), .B(N460), .C(
        N459), .Y(ADD_26x26_fast_I210_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I71_Y (.A(N324), .B(N321), .Y(
        N439));
    DFN1E0C0 \integ[20]  (.D(\un1_integ[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[20]_net_1 ));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I244_Y (.A(\state_0[0]_net_1 ), 
        .B(LED_5[7]), .C(N640), .Y(\un1_integ[14] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I207_Y_1 (.A(N404), .B(N400), .C(
        N461), .Y(ADD_26x26_fast_I207_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I106_Y (.A(N428), .B(N425), .C(
        N424), .Y(N477));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_1 (.A(
        ADD_26x26_fast_I208_un1_Y_0), .B(N541), .C(
        ADD_26x26_fast_I208_Y_0), .Y(ADD_26x26_fast_I208_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I102_Y (.A(N424), .B(N421), .C(
        N420), .Y(N473));
    AX1D un1_integ_0_0_ADD_26x26_fast_I251_Y (.A(I176_un1_Y), .B(
        ADD_26x26_fast_I208_Y_1), .C(ADD_26x26_fast_I251_Y_0), .Y(
        \un1_integ[21] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I121_un1_Y (.A(N441), .B(
        \state_RNI74E11[0]_net_1 ), .Y(I121_un1_Y));
    DFN1E0C0 \integ[18]  (.D(\un1_integ[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[18]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I4_P0N (.A(average[4]), .B(
        \state_RNIFCE11[0]_net_1 ), .Y(N330));
    AO1 un1_integ_0_0_ADD_26x26_fast_I144_Y (.A(N468), .B(N475), .C(
        N467), .Y(N521));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_0 (.A(N465), .B(N458), .C(
        N457), .Y(ADD_26x26_fast_I209_Y_0));
    NOR2A \state_RNIRF3H[1]  (.A(\state[1]_net_1 ), .B(avg_old[5]), .Y(
        \un18_next_int_m[5] ));
    OR2 \state_RNIB8E11[0]  (.A(\inf_abs0_m[2] ), .B(
        \un18_next_int_m[2] ), .Y(\state_RNIB8E11[0]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I148_Y (.A(I148_un1_Y), .B(N471), 
        .Y(N525));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I60_Y (.A(N335), .B(
        \state_RNILIE11[0]_net_1 ), .C(LED_5[0]), .Y(N428));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y (.A(
        ADD_26x26_fast_I232_Y_0), .B(N493), .Y(\un1_integ[2] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I204_Y_2 (.A(N398), .B(
        ADD_26x26_fast_I204_Y_0), .C(N455), .Y(ADD_26x26_fast_I204_Y_2)
        );
    DFN1C0 \state[1]  (.D(\state_RNO_5[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[1]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I110_un1_Y (.A(N432), .B(N429), 
        .Y(I110_un1_Y));
    OA1 un1_integ_0_0_ADD_26x26_fast_I9_G0N (.A(\un18_next_int_m[9] ), 
        .B(\inf_abs0_m[9] ), .C(LED_5[2]), .Y(N344));
    OA1B un1_integ_0_0_ADD_26x26_fast_I40_Y (.A(\integ[17]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N408));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I65_Y (.A(N333), .B(N330), .Y(
        N433));
    NOR2A \state_RNINB3H[1]  (.A(\state[1]_net_1 ), .B(avg_old[1]), .Y(
        \un18_next_int_m[1] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I188_Y (.A(N522), .B(N537), .C(
        N521), .Y(N637));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I178_un1_Y (.A(N512), .B(N527), 
        .Y(I178_un1_Y));
    AO1B un1_integ_0_0_ADD_26x26_fast_I45_Y (.A(LED_5[7]), .B(
        \integ[15]_net_1 ), .C(\state_1[0]_net_1 ), .Y(N413));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I137_Y (.A(N468), .B(N460), .Y(
        N514));
    OR2 un1_integ_0_0_ADD_26x26_fast_I3_P0N (.A(average[3]), .B(
        \un1_next_int[3] ), .Y(N327));
    OR2 \state_RNIJGE11[0]  (.A(\un18_next_int_m[6] ), .B(
        \inf_abs0_m[6] ), .Y(\un1_next_int[6] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I50_Y (.A(N350), .B(N354), .C(
        N353), .Y(N418));
    AO1 un1_integ_0_0_ADD_26x26_fast_I204_Y_3 (.A(N517), .B(N502), .C(
        ADD_26x26_fast_I204_Y_2), .Y(ADD_26x26_fast_I204_Y_3));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I74_un1_Y (.A(N318), .B(
        \state_RNI74E11[0]_net_1 ), .Y(I74_un1_Y));
    OA1B un1_integ_0_0_ADD_26x26_fast_I36_Y (.A(\integ[18]_net_1 ), .B(
        \integ[19]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N404));
    NOR2B \state_RNIMUAG[0]  (.A(avg_new[5]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[5] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I0_P0N (.A(\integ[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(N318));
    OR2 \state_RNIHEE11[0]  (.A(\un18_next_int_m[5] ), .B(
        \inf_abs0_m[5] ), .Y(\un1_next_int[5] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I55_Y (.A(N348), .B(N345), .Y(
        N423));
    OA1 un1_integ_0_0_ADD_26x26_fast_I205_un1_Y (.A(N535), .B(
        I195_un1_Y), .C(ADD_26x26_fast_I205_un1_Y_0), .Y(I205_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I163_un1_Y (.A(N490), .B(
        \state_RNI74E11[0]_net_1 ), .Y(I163_un1_Y));
    NOR2B \state_1_RNIIA8G[0]  (.A(avg_new[10]), .B(\state_1[0]_net_1 )
        , .Y(\inf_abs0_m[10] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I206_Y_1 (.A(N402), .B(N398), .C(
        N459), .Y(ADD_26x26_fast_I206_Y_1));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I5_G0N (.A(average[5]), .B(
        \un1_next_int[5] ), .Y(N332));
    DFN1E0C0 \integ[7]  (.D(\un1_integ[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(LED_5[0]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_2 (.A(N508), .B(N523), .C(
        ADD_26x26_fast_I207_Y_1), .Y(ADD_26x26_fast_I207_Y_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I4_G0N (.A(average[4]), .B(
        \state_RNIFCE11[0]_net_1 ), .Y(N329));
    OR2 \state_RNIRSHK[1]  (.A(\un18_next_int_m[11] ), .B(
        \inf_abs0_m[11] ), .Y(\un1_next_int[11] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y (.A(
        ADD_26x26_fast_I234_Y_0), .B(N543), .Y(\un1_integ[4] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I205_Y_2 (.A(
        ADD_26x26_fast_I205_Y_1), .B(N457), .Y(ADD_26x26_fast_I205_Y_2)
        );
    NOR2B un1_integ_0_0_ADD_26x26_fast_I162_un1_Y (.A(N488), .B(N442), 
        .Y(I162_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I240_Y (.A(N531), .B(I193_un1_Y), 
        .C(ADD_26x26_fast_I240_Y_0), .Y(\un1_integ[10] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I156_Y (.A(N487), .B(N480), .C(
        N479), .Y(N533));
    DFN1E0C0 \integ[8]  (.D(\un1_integ[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(LED_5[1]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I85_Y (.A(N403), .B(N407), .Y(
        N456));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I251_Y_0 (.A(\integ[21]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I251_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I152_Y (.A(I152_un1_Y), .B(N475), 
        .Y(N529));
    OR3 un1_integ_0_0_ADD_26x26_fast_I9_P0N (.A(\un18_next_int_m[9] ), 
        .B(\inf_abs0_m[9] ), .C(LED_5[2]), .Y(N345));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I208_un1_Y_0 (.A(N510), .B(N526)
        , .Y(ADD_26x26_fast_I208_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I191_Y (.A(N528), .B(N543), .C(
        N527), .Y(N646));
    AO1B un1_integ_0_0_ADD_26x26_fast_I31_Y (.A(\integ[21]_net_1 ), .B(
        \integ[22]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N399));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I206_un1_Y (.A(N522), .B(N506), 
        .C(N537), .Y(I206_un1_Y));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I235_Y_0 (.A(average[5]), .B(
        \un1_next_int[5] ), .Y(ADD_26x26_fast_I235_Y_0));
    NOR2A \state_RNIQE3H[1]  (.A(\state[1]_net_1 ), .B(avg_old[4]), .Y(
        \un18_next_int_m[4] ));
    NOR2 \state_0_RNISJ4B[0]  (.A(\state[1]_net_1 ), .B(
        \state_0[0]_net_1 ), .Y(avg_done_0));
    NOR2B \state_RNIHPAG[0]  (.A(avg_new[0]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[0] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I241_Y (.A(N529), .B(I192_un1_Y), 
        .C(ADD_26x26_fast_I241_Y_0), .Y(\un1_integ[11] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I11_P0N (.A(\un1_next_int[11] ), 
        .B(LED_5[4]), .Y(N351));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I105_Y (.A(N423), .B(N427), .Y(
        N476));
    AO1 un1_integ_0_0_ADD_26x26_fast_I213_Y_0 (.A(
        ADD_26x26_fast_I213_un1_Y_0), .B(N520), .C(N519), .Y(
        ADD_26x26_fast_I213_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I238_Y_0 (.A(LED_5[1]), .B(
        \un1_next_int[8] ), .Y(ADD_26x26_fast_I238_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I101_Y (.A(N423), .B(N419), .Y(
        N472));
    NOR2A \state_RNI7G94[1]  (.A(\state[1]_net_1 ), .B(avg_old[10]), 
        .Y(\un18_next_int_m[10] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I66_Y (.A(N326), .B(N330), .C(
        N329), .Y(N434));
    AX1D un1_integ_0_0_ADD_26x26_fast_I248_Y (.A(I182_un1_Y), .B(
        ADD_26x26_fast_I211_Y_1), .C(ADD_26x26_fast_I248_Y_0), .Y(
        \un1_integ[18] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I99_Y (.A(N417), .B(N421), .Y(
        N470));
    AO1 un1_integ_0_0_ADD_26x26_fast_I92_Y (.A(N411), .B(N414), .C(
        N410), .Y(N463));
    AO1 un1_integ_0_0_ADD_26x26_fast_I72_Y (.A(N317), .B(N321), .C(
        N320), .Y(N440));
    OR2A un1_integ_0_0_ADD_26x26_fast_I13_P0N (.A(\state_1[0]_net_1 ), 
        .B(LED_5[6]), .Y(N357));
    OA1B un1_integ_0_0_ADD_26x26_fast_I46_Y (.A(LED_5[7]), .B(LED_5[6])
        , .C(\state_1[0]_net_1 ), .Y(N414));
    NOR2B \state_1_RNIQNJE[0]  (.A(avg_done), .B(calc_avg), .Y(
        \state_1_RNIQNJE[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I116_Y (.A(N438), .B(N435), .C(
        N434), .Y(N487));
    OR2 un1_integ_0_0_ADD_26x26_fast_I112_Y (.A(I112_un1_Y), .B(N430), 
        .Y(N483));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I8_G0N (.A(\un1_next_int[8] ), 
        .B(LED_5[1]), .Y(N341));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I213_un1_Y_0 (.A(N482), .B(N490)
        , .C(\state_RNI74E11[0]_net_1 ), .Y(
        ADD_26x26_fast_I213_un1_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y_0 (.A(average[4]), .B(
        \state_RNIFCE11[0]_net_1 ), .Y(ADD_26x26_fast_I234_Y_0));
    
endmodule


module error_sr_13s_5s_2(
       cur_vd,
       avg_new,
       avg_old,
       avg_enable_1,
       avg_enable_0,
       avg_enable,
       n_rst_c,
       clk_c
    );
input  [11:0] cur_vd;
output [11:0] avg_new;
output [11:0] avg_old;
input  avg_enable_1;
input  avg_enable_0;
input  avg_enable;
input  n_rst_c;
input  clk_c;

    wire \sr_3_[0]_net_1 , \sr_3_[1]_net_1 , \sr_3_[2]_net_1 , 
        \sr_3_[3]_net_1 , \sr_3_[4]_net_1 , \sr_3_[5]_net_1 , 
        \sr_3_[6]_net_1 , \sr_3_[7]_net_1 , \sr_3_[8]_net_1 , 
        \sr_3_[9]_net_1 , \sr_3_[10]_net_1 , \sr_3_[11]_net_1 , 
        \sr_2_[0]_net_1 , \sr_2_[1]_net_1 , \sr_2_[2]_net_1 , 
        \sr_2_[3]_net_1 , \sr_2_[4]_net_1 , \sr_2_[5]_net_1 , 
        \sr_2_[6]_net_1 , \sr_2_[7]_net_1 , \sr_2_[8]_net_1 , 
        \sr_2_[9]_net_1 , \sr_2_[10]_net_1 , \sr_2_[11]_net_1 , 
        \sr_1_[0]_net_1 , \sr_1_[1]_net_1 , \sr_1_[2]_net_1 , 
        \sr_1_[3]_net_1 , \sr_1_[4]_net_1 , \sr_1_[5]_net_1 , 
        \sr_1_[6]_net_1 , \sr_1_[7]_net_1 , \sr_1_[8]_net_1 , 
        \sr_1_[9]_net_1 , \sr_1_[10]_net_1 , \sr_1_[11]_net_1 , GND, 
        VCC;
    
    DFN1E1C0 \sr_1_[11]  (.D(avg_new[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[11]_net_1 ));
    DFN1E1C0 \sr_3_[3]  (.D(\sr_2_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[3]_net_1 ));
    DFN1E1C0 \sr_4_[4]  (.D(\sr_3_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[4]));
    DFN1E1C0 \sr_0_[10]  (.D(cur_vd[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(avg_new[10]));
    DFN1E1C0 \sr_4_[8]  (.D(\sr_3_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[8]));
    DFN1E1C0 \sr_4_[0]  (.D(\sr_3_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[0]));
    DFN1E1C0 \sr_1_[2]  (.D(avg_new[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[2]_net_1 ));
    DFN1E1C0 \sr_0_[2]  (.D(cur_vd[2]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[2]));
    DFN1E1C0 \sr_2_[2]  (.D(\sr_1_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[2]_net_1 ));
    DFN1E1C0 \sr_0_[11]  (.D(cur_vd[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(avg_new[11]));
    DFN1E1C0 \sr_1_[3]  (.D(avg_new[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[3]_net_1 ));
    DFN1E1C0 \sr_0_[3]  (.D(cur_vd[3]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[3]));
    DFN1E1C0 \sr_1_[10]  (.D(avg_new[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[10]_net_1 ));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \sr_4_[10]  (.D(\sr_3_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[10]));
    DFN1E1C0 \sr_3_[11]  (.D(\sr_2_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[11]_net_1 ));
    DFN1E1C0 \sr_2_[3]  (.D(\sr_1_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[3]_net_1 ));
    DFN1E1C0 \sr_3_[6]  (.D(\sr_2_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[6]_net_1 ));
    DFN1E1C0 \sr_3_[1]  (.D(\sr_2_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[1]_net_1 ));
    DFN1E1C0 \sr_4_[2]  (.D(\sr_3_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[2]));
    DFN1E1C0 \sr_1_[6]  (.D(avg_new[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[6]_net_1 ));
    DFN1E1C0 \sr_4_[3]  (.D(\sr_3_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[3]));
    DFN1E1C0 \sr_0_[6]  (.D(cur_vd[6]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[6]));
    DFN1E1C0 \sr_3_[9]  (.D(\sr_2_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[9]_net_1 ));
    DFN1E1C0 \sr_1_[1]  (.D(avg_new[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[1]_net_1 ));
    DFN1E1C0 \sr_0_[1]  (.D(cur_vd[1]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[1]));
    DFN1E1C0 \sr_2_[6]  (.D(\sr_1_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[6]_net_1 ));
    DFN1E1C0 \sr_2_[1]  (.D(\sr_1_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[1]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1C0 \sr_3_[5]  (.D(\sr_2_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[5]_net_1 ));
    DFN1E1C0 \sr_3_[7]  (.D(\sr_2_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[7]_net_1 ));
    DFN1E1C0 \sr_1_[9]  (.D(avg_new[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[9]_net_1 ));
    DFN1E1C0 \sr_0_[9]  (.D(cur_vd[9]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[9]));
    DFN1E1C0 \sr_2_[11]  (.D(\sr_1_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[11]_net_1 ));
    DFN1E1C0 \sr_4_[6]  (.D(\sr_3_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[6]));
    DFN1E1C0 \sr_2_[9]  (.D(\sr_1_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[9]_net_1 ));
    DFN1E1C0 \sr_4_[11]  (.D(\sr_3_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[11]));
    DFN1E1C0 \sr_4_[1]  (.D(\sr_3_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[1]));
    DFN1E1C0 \sr_3_[4]  (.D(\sr_2_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[4]_net_1 ));
    DFN1E1C0 \sr_1_[5]  (.D(avg_new[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[5]_net_1 ));
    DFN1E1C0 \sr_0_[5]  (.D(cur_vd[5]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[5]));
    DFN1E1C0 \sr_1_[7]  (.D(avg_new[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[7]_net_1 ));
    DFN1E1C0 \sr_0_[7]  (.D(cur_vd[7]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[7]));
    DFN1E1C0 \sr_3_[8]  (.D(\sr_2_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[8]_net_1 ));
    DFN1E1C0 \sr_3_[0]  (.D(\sr_2_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[0]_net_1 ));
    DFN1E1C0 \sr_2_[5]  (.D(\sr_1_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[5]_net_1 ));
    DFN1E1C0 \sr_2_[7]  (.D(\sr_1_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[7]_net_1 ));
    DFN1E1C0 \sr_4_[9]  (.D(\sr_3_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[9]));
    DFN1E1C0 \sr_1_[4]  (.D(avg_new[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[4]_net_1 ));
    DFN1E1C0 \sr_0_[4]  (.D(cur_vd[4]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[4]));
    DFN1E1C0 \sr_1_[8]  (.D(avg_new[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[8]_net_1 ));
    DFN1E1C0 \sr_1_[0]  (.D(avg_new[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[0]_net_1 ));
    DFN1E1C0 \sr_2_[4]  (.D(\sr_1_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[4]_net_1 ));
    DFN1E1C0 \sr_0_[8]  (.D(cur_vd[8]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[8]));
    DFN1E1C0 \sr_0_[0]  (.D(cur_vd[0]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[0]));
    DFN1E1C0 \sr_4_[5]  (.D(\sr_3_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[5]));
    DFN1E1C0 \sr_2_[8]  (.D(\sr_1_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[8]_net_1 ));
    DFN1E1C0 \sr_2_[0]  (.D(\sr_1_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[0]_net_1 ));
    DFN1E1C0 \sr_4_[7]  (.D(\sr_3_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[7]));
    DFN1E1C0 \sr_3_[10]  (.D(\sr_2_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[10]_net_1 ));
    DFN1E1C0 \sr_3_[2]  (.D(\sr_2_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[2]_net_1 ));
    DFN1E1C0 \sr_2_[10]  (.D(\sr_1_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[10]_net_1 ));
    
endmodule


module error_sr_13s_64s_2(
       sr_old,
       sr_new,
       cur_error,
       sr_prev,
       sr_new_0_0,
       sr_new_1_0,
       int_enable,
       n_rst_c,
       clk_c
    );
output [12:0] sr_old;
output [12:0] sr_new;
input  [12:0] cur_error;
output [12:0] sr_prev;
output sr_new_0_0;
output sr_new_1_0;
input  int_enable;
input  n_rst_c;
input  clk_c;

    wire \sr_9_[0]_net_1 , \sr_8_[0]_net_1 , \sr_9_[1]_net_1 , 
        \sr_8_[1]_net_1 , \sr_9_[2]_net_1 , \sr_8_[2]_net_1 , 
        \sr_9_[3]_net_1 , \sr_8_[3]_net_1 , \sr_9_[4]_net_1 , 
        \sr_8_[4]_net_1 , \sr_9_[5]_net_1 , \sr_8_[5]_net_1 , 
        \sr_9_[6]_net_1 , \sr_8_[6]_net_1 , \sr_9_[7]_net_1 , 
        \sr_8_[7]_net_1 , \sr_9_[8]_net_1 , \sr_8_[8]_net_1 , 
        \sr_9_[9]_net_1 , \sr_8_[9]_net_1 , \sr_9_[10]_net_1 , 
        \sr_8_[10]_net_1 , \sr_9_[11]_net_1 , \sr_8_[11]_net_1 , 
        \sr_9_[12]_net_1 , \sr_8_[12]_net_1 , \sr_7_[0]_net_1 , 
        \sr_7_[1]_net_1 , \sr_7_[2]_net_1 , \sr_7_[3]_net_1 , 
        \sr_7_[4]_net_1 , \sr_7_[5]_net_1 , \sr_7_[6]_net_1 , 
        \sr_7_[7]_net_1 , \sr_7_[8]_net_1 , \sr_7_[9]_net_1 , 
        \sr_7_[10]_net_1 , \sr_7_[11]_net_1 , \sr_7_[12]_net_1 , 
        \sr_6_[0]_net_1 , \sr_6_[1]_net_1 , \sr_6_[2]_net_1 , 
        \sr_6_[3]_net_1 , \sr_6_[4]_net_1 , \sr_6_[5]_net_1 , 
        \sr_6_[6]_net_1 , \sr_6_[7]_net_1 , \sr_6_[8]_net_1 , 
        \sr_6_[9]_net_1 , \sr_6_[10]_net_1 , \sr_6_[11]_net_1 , 
        \sr_6_[12]_net_1 , \sr_5_[0]_net_1 , \sr_5_[1]_net_1 , 
        \sr_5_[2]_net_1 , \sr_5_[3]_net_1 , \sr_5_[4]_net_1 , 
        \sr_5_[5]_net_1 , \sr_5_[6]_net_1 , \sr_5_[7]_net_1 , 
        \sr_5_[8]_net_1 , \sr_5_[9]_net_1 , \sr_5_[10]_net_1 , 
        \sr_5_[11]_net_1 , \sr_5_[12]_net_1 , \sr_4_[0]_net_1 , 
        \sr_4_[1]_net_1 , \sr_4_[2]_net_1 , \sr_4_[3]_net_1 , 
        \sr_4_[4]_net_1 , \sr_4_[5]_net_1 , \sr_4_[6]_net_1 , 
        \sr_4_[7]_net_1 , \sr_4_[8]_net_1 , \sr_4_[9]_net_1 , 
        \sr_4_[10]_net_1 , \sr_4_[11]_net_1 , \sr_4_[12]_net_1 , 
        \sr_3_[0]_net_1 , \sr_3_[1]_net_1 , \sr_3_[2]_net_1 , 
        \sr_3_[3]_net_1 , \sr_3_[4]_net_1 , \sr_3_[5]_net_1 , 
        \sr_3_[6]_net_1 , \sr_3_[7]_net_1 , \sr_3_[8]_net_1 , 
        \sr_3_[9]_net_1 , \sr_3_[10]_net_1 , \sr_3_[11]_net_1 , 
        \sr_3_[12]_net_1 , \sr_2_[0]_net_1 , \sr_2_[1]_net_1 , 
        \sr_2_[2]_net_1 , \sr_2_[3]_net_1 , \sr_2_[4]_net_1 , 
        \sr_2_[5]_net_1 , \sr_2_[6]_net_1 , \sr_2_[7]_net_1 , 
        \sr_2_[8]_net_1 , \sr_2_[9]_net_1 , \sr_2_[10]_net_1 , 
        \sr_2_[11]_net_1 , \sr_2_[12]_net_1 , \sr_24_[0]_net_1 , 
        \sr_23_[0]_net_1 , \sr_24_[1]_net_1 , \sr_23_[1]_net_1 , 
        \sr_24_[2]_net_1 , \sr_23_[2]_net_1 , \sr_24_[3]_net_1 , 
        \sr_23_[3]_net_1 , \sr_24_[4]_net_1 , \sr_23_[4]_net_1 , 
        \sr_24_[5]_net_1 , \sr_23_[5]_net_1 , \sr_24_[6]_net_1 , 
        \sr_23_[6]_net_1 , \sr_24_[7]_net_1 , \sr_23_[7]_net_1 , 
        \sr_24_[8]_net_1 , \sr_23_[8]_net_1 , \sr_24_[9]_net_1 , 
        \sr_23_[9]_net_1 , \sr_24_[10]_net_1 , \sr_23_[10]_net_1 , 
        \sr_24_[11]_net_1 , \sr_23_[11]_net_1 , \sr_24_[12]_net_1 , 
        \sr_23_[12]_net_1 , \sr_22_[0]_net_1 , \sr_22_[1]_net_1 , 
        \sr_22_[2]_net_1 , \sr_22_[3]_net_1 , \sr_22_[4]_net_1 , 
        \sr_22_[5]_net_1 , \sr_22_[6]_net_1 , \sr_22_[7]_net_1 , 
        \sr_22_[8]_net_1 , \sr_22_[9]_net_1 , \sr_22_[10]_net_1 , 
        \sr_22_[11]_net_1 , \sr_22_[12]_net_1 , \sr_21_[0]_net_1 , 
        \sr_21_[1]_net_1 , \sr_21_[2]_net_1 , \sr_21_[3]_net_1 , 
        \sr_21_[4]_net_1 , \sr_21_[5]_net_1 , \sr_21_[6]_net_1 , 
        \sr_21_[7]_net_1 , \sr_21_[8]_net_1 , \sr_21_[9]_net_1 , 
        \sr_21_[10]_net_1 , \sr_21_[11]_net_1 , \sr_21_[12]_net_1 , 
        \sr_20_[0]_net_1 , \sr_20_[1]_net_1 , \sr_20_[2]_net_1 , 
        \sr_20_[3]_net_1 , \sr_20_[4]_net_1 , \sr_20_[5]_net_1 , 
        \sr_20_[6]_net_1 , \sr_20_[7]_net_1 , \sr_20_[8]_net_1 , 
        \sr_20_[9]_net_1 , \sr_20_[10]_net_1 , \sr_20_[11]_net_1 , 
        \sr_20_[12]_net_1 , \sr_19_[0]_net_1 , \sr_19_[1]_net_1 , 
        \sr_19_[2]_net_1 , \sr_19_[3]_net_1 , \sr_19_[4]_net_1 , 
        \sr_19_[5]_net_1 , \sr_19_[6]_net_1 , \sr_19_[7]_net_1 , 
        \sr_19_[8]_net_1 , \sr_19_[9]_net_1 , \sr_19_[10]_net_1 , 
        \sr_19_[11]_net_1 , \sr_19_[12]_net_1 , \sr_18_[0]_net_1 , 
        \sr_18_[1]_net_1 , \sr_18_[2]_net_1 , \sr_18_[3]_net_1 , 
        \sr_18_[4]_net_1 , \sr_18_[5]_net_1 , \sr_18_[6]_net_1 , 
        \sr_18_[7]_net_1 , \sr_18_[8]_net_1 , \sr_18_[9]_net_1 , 
        \sr_18_[10]_net_1 , \sr_18_[11]_net_1 , \sr_18_[12]_net_1 , 
        \sr_17_[0]_net_1 , \sr_17_[1]_net_1 , \sr_17_[2]_net_1 , 
        \sr_17_[3]_net_1 , \sr_17_[4]_net_1 , \sr_17_[5]_net_1 , 
        \sr_17_[6]_net_1 , \sr_17_[7]_net_1 , \sr_17_[8]_net_1 , 
        \sr_17_[9]_net_1 , \sr_17_[10]_net_1 , \sr_17_[11]_net_1 , 
        \sr_17_[12]_net_1 , \sr_16_[0]_net_1 , \sr_16_[1]_net_1 , 
        \sr_16_[2]_net_1 , \sr_16_[3]_net_1 , \sr_16_[4]_net_1 , 
        \sr_16_[5]_net_1 , \sr_16_[6]_net_1 , \sr_16_[7]_net_1 , 
        \sr_16_[8]_net_1 , \sr_16_[9]_net_1 , \sr_16_[10]_net_1 , 
        \sr_16_[11]_net_1 , \sr_16_[12]_net_1 , \sr_15_[0]_net_1 , 
        \sr_15_[1]_net_1 , \sr_15_[2]_net_1 , \sr_15_[3]_net_1 , 
        \sr_15_[4]_net_1 , \sr_15_[5]_net_1 , \sr_15_[6]_net_1 , 
        \sr_15_[7]_net_1 , \sr_15_[8]_net_1 , \sr_15_[9]_net_1 , 
        \sr_15_[10]_net_1 , \sr_15_[11]_net_1 , \sr_15_[12]_net_1 , 
        \sr_14_[0]_net_1 , \sr_14_[1]_net_1 , \sr_14_[2]_net_1 , 
        \sr_14_[3]_net_1 , \sr_14_[4]_net_1 , \sr_14_[5]_net_1 , 
        \sr_14_[6]_net_1 , \sr_14_[7]_net_1 , \sr_14_[8]_net_1 , 
        \sr_14_[9]_net_1 , \sr_14_[10]_net_1 , \sr_14_[11]_net_1 , 
        \sr_14_[12]_net_1 , \sr_13_[0]_net_1 , \sr_13_[1]_net_1 , 
        \sr_13_[2]_net_1 , \sr_13_[3]_net_1 , \sr_13_[4]_net_1 , 
        \sr_13_[5]_net_1 , \sr_13_[6]_net_1 , \sr_13_[7]_net_1 , 
        \sr_13_[8]_net_1 , \sr_13_[9]_net_1 , \sr_13_[10]_net_1 , 
        \sr_13_[11]_net_1 , \sr_13_[12]_net_1 , \sr_12_[0]_net_1 , 
        \sr_12_[1]_net_1 , \sr_12_[2]_net_1 , \sr_12_[3]_net_1 , 
        \sr_12_[4]_net_1 , \sr_12_[5]_net_1 , \sr_12_[6]_net_1 , 
        \sr_12_[7]_net_1 , \sr_12_[8]_net_1 , \sr_12_[9]_net_1 , 
        \sr_12_[10]_net_1 , \sr_12_[11]_net_1 , \sr_12_[12]_net_1 , 
        \sr_11_[0]_net_1 , \sr_11_[1]_net_1 , \sr_11_[2]_net_1 , 
        \sr_11_[3]_net_1 , \sr_11_[4]_net_1 , \sr_11_[5]_net_1 , 
        \sr_11_[6]_net_1 , \sr_11_[7]_net_1 , \sr_11_[8]_net_1 , 
        \sr_11_[9]_net_1 , \sr_11_[10]_net_1 , \sr_11_[11]_net_1 , 
        \sr_11_[12]_net_1 , \sr_10_[0]_net_1 , \sr_10_[1]_net_1 , 
        \sr_10_[2]_net_1 , \sr_10_[3]_net_1 , \sr_10_[4]_net_1 , 
        \sr_10_[5]_net_1 , \sr_10_[6]_net_1 , \sr_10_[7]_net_1 , 
        \sr_10_[8]_net_1 , \sr_10_[9]_net_1 , \sr_10_[10]_net_1 , 
        \sr_10_[11]_net_1 , \sr_10_[12]_net_1 , \sr_39_[0]_net_1 , 
        \sr_38_[0]_net_1 , \sr_39_[1]_net_1 , \sr_38_[1]_net_1 , 
        \sr_39_[2]_net_1 , \sr_38_[2]_net_1 , \sr_39_[3]_net_1 , 
        \sr_38_[3]_net_1 , \sr_39_[4]_net_1 , \sr_38_[4]_net_1 , 
        \sr_39_[5]_net_1 , \sr_38_[5]_net_1 , \sr_39_[6]_net_1 , 
        \sr_38_[6]_net_1 , \sr_39_[7]_net_1 , \sr_38_[7]_net_1 , 
        \sr_39_[8]_net_1 , \sr_38_[8]_net_1 , \sr_39_[9]_net_1 , 
        \sr_38_[9]_net_1 , \sr_39_[10]_net_1 , \sr_38_[10]_net_1 , 
        \sr_39_[11]_net_1 , \sr_38_[11]_net_1 , \sr_39_[12]_net_1 , 
        \sr_38_[12]_net_1 , \sr_37_[0]_net_1 , \sr_37_[1]_net_1 , 
        \sr_37_[2]_net_1 , \sr_37_[3]_net_1 , \sr_37_[4]_net_1 , 
        \sr_37_[5]_net_1 , \sr_37_[6]_net_1 , \sr_37_[7]_net_1 , 
        \sr_37_[8]_net_1 , \sr_37_[9]_net_1 , \sr_37_[10]_net_1 , 
        \sr_37_[11]_net_1 , \sr_37_[12]_net_1 , \sr_36_[0]_net_1 , 
        \sr_36_[1]_net_1 , \sr_36_[2]_net_1 , \sr_36_[3]_net_1 , 
        \sr_36_[4]_net_1 , \sr_36_[5]_net_1 , \sr_36_[6]_net_1 , 
        \sr_36_[7]_net_1 , \sr_36_[8]_net_1 , \sr_36_[9]_net_1 , 
        \sr_36_[10]_net_1 , \sr_36_[11]_net_1 , \sr_36_[12]_net_1 , 
        \sr_35_[0]_net_1 , \sr_35_[1]_net_1 , \sr_35_[2]_net_1 , 
        \sr_35_[3]_net_1 , \sr_35_[4]_net_1 , \sr_35_[5]_net_1 , 
        \sr_35_[6]_net_1 , \sr_35_[7]_net_1 , \sr_35_[8]_net_1 , 
        \sr_35_[9]_net_1 , \sr_35_[10]_net_1 , \sr_35_[11]_net_1 , 
        \sr_35_[12]_net_1 , \sr_34_[0]_net_1 , \sr_34_[1]_net_1 , 
        \sr_34_[2]_net_1 , \sr_34_[3]_net_1 , \sr_34_[4]_net_1 , 
        \sr_34_[5]_net_1 , \sr_34_[6]_net_1 , \sr_34_[7]_net_1 , 
        \sr_34_[8]_net_1 , \sr_34_[9]_net_1 , \sr_34_[10]_net_1 , 
        \sr_34_[11]_net_1 , \sr_34_[12]_net_1 , \sr_33_[0]_net_1 , 
        \sr_33_[1]_net_1 , \sr_33_[2]_net_1 , \sr_33_[3]_net_1 , 
        \sr_33_[4]_net_1 , \sr_33_[5]_net_1 , \sr_33_[6]_net_1 , 
        \sr_33_[7]_net_1 , \sr_33_[8]_net_1 , \sr_33_[9]_net_1 , 
        \sr_33_[10]_net_1 , \sr_33_[11]_net_1 , \sr_33_[12]_net_1 , 
        \sr_32_[0]_net_1 , \sr_32_[1]_net_1 , \sr_32_[2]_net_1 , 
        \sr_32_[3]_net_1 , \sr_32_[4]_net_1 , \sr_32_[5]_net_1 , 
        \sr_32_[6]_net_1 , \sr_32_[7]_net_1 , \sr_32_[8]_net_1 , 
        \sr_32_[9]_net_1 , \sr_32_[10]_net_1 , \sr_32_[11]_net_1 , 
        \sr_32_[12]_net_1 , \sr_31_[0]_net_1 , \sr_31_[1]_net_1 , 
        \sr_31_[2]_net_1 , \sr_31_[3]_net_1 , \sr_31_[4]_net_1 , 
        \sr_31_[5]_net_1 , \sr_31_[6]_net_1 , \sr_31_[7]_net_1 , 
        \sr_31_[8]_net_1 , \sr_31_[9]_net_1 , \sr_31_[10]_net_1 , 
        \sr_31_[11]_net_1 , \sr_31_[12]_net_1 , \sr_30_[0]_net_1 , 
        \sr_30_[1]_net_1 , \sr_30_[2]_net_1 , \sr_30_[3]_net_1 , 
        \sr_30_[4]_net_1 , \sr_30_[5]_net_1 , \sr_30_[6]_net_1 , 
        \sr_30_[7]_net_1 , \sr_30_[8]_net_1 , \sr_30_[9]_net_1 , 
        \sr_30_[10]_net_1 , \sr_30_[11]_net_1 , \sr_30_[12]_net_1 , 
        \sr_29_[0]_net_1 , \sr_29_[1]_net_1 , \sr_29_[2]_net_1 , 
        \sr_29_[3]_net_1 , \sr_29_[4]_net_1 , \sr_29_[5]_net_1 , 
        \sr_29_[6]_net_1 , \sr_29_[7]_net_1 , \sr_29_[8]_net_1 , 
        \sr_29_[9]_net_1 , \sr_29_[10]_net_1 , \sr_29_[11]_net_1 , 
        \sr_29_[12]_net_1 , \sr_28_[0]_net_1 , \sr_28_[1]_net_1 , 
        \sr_28_[2]_net_1 , \sr_28_[3]_net_1 , \sr_28_[4]_net_1 , 
        \sr_28_[5]_net_1 , \sr_28_[6]_net_1 , \sr_28_[7]_net_1 , 
        \sr_28_[8]_net_1 , \sr_28_[9]_net_1 , \sr_28_[10]_net_1 , 
        \sr_28_[11]_net_1 , \sr_28_[12]_net_1 , \sr_27_[0]_net_1 , 
        \sr_27_[1]_net_1 , \sr_27_[2]_net_1 , \sr_27_[3]_net_1 , 
        \sr_27_[4]_net_1 , \sr_27_[5]_net_1 , \sr_27_[6]_net_1 , 
        \sr_27_[7]_net_1 , \sr_27_[8]_net_1 , \sr_27_[9]_net_1 , 
        \sr_27_[10]_net_1 , \sr_27_[11]_net_1 , \sr_27_[12]_net_1 , 
        \sr_26_[0]_net_1 , \sr_26_[1]_net_1 , \sr_26_[2]_net_1 , 
        \sr_26_[3]_net_1 , \sr_26_[4]_net_1 , \sr_26_[5]_net_1 , 
        \sr_26_[6]_net_1 , \sr_26_[7]_net_1 , \sr_26_[8]_net_1 , 
        \sr_26_[9]_net_1 , \sr_26_[10]_net_1 , \sr_26_[11]_net_1 , 
        \sr_26_[12]_net_1 , \sr_25_[0]_net_1 , \sr_25_[1]_net_1 , 
        \sr_25_[2]_net_1 , \sr_25_[3]_net_1 , \sr_25_[4]_net_1 , 
        \sr_25_[5]_net_1 , \sr_25_[6]_net_1 , \sr_25_[7]_net_1 , 
        \sr_25_[8]_net_1 , \sr_25_[9]_net_1 , \sr_25_[10]_net_1 , 
        \sr_25_[11]_net_1 , \sr_25_[12]_net_1 , \sr_54_[0]_net_1 , 
        \sr_53_[0]_net_1 , \sr_54_[1]_net_1 , \sr_53_[1]_net_1 , 
        \sr_54_[2]_net_1 , \sr_53_[2]_net_1 , \sr_54_[3]_net_1 , 
        \sr_53_[3]_net_1 , \sr_54_[4]_net_1 , \sr_53_[4]_net_1 , 
        \sr_54_[5]_net_1 , \sr_53_[5]_net_1 , \sr_54_[6]_net_1 , 
        \sr_53_[6]_net_1 , \sr_54_[7]_net_1 , \sr_53_[7]_net_1 , 
        \sr_54_[8]_net_1 , \sr_53_[8]_net_1 , \sr_54_[9]_net_1 , 
        \sr_53_[9]_net_1 , \sr_54_[10]_net_1 , \sr_53_[10]_net_1 , 
        \sr_54_[11]_net_1 , \sr_53_[11]_net_1 , \sr_54_[12]_net_1 , 
        \sr_53_[12]_net_1 , \sr_52_[0]_net_1 , \sr_52_[1]_net_1 , 
        \sr_52_[2]_net_1 , \sr_52_[3]_net_1 , \sr_52_[4]_net_1 , 
        \sr_52_[5]_net_1 , \sr_52_[6]_net_1 , \sr_52_[7]_net_1 , 
        \sr_52_[8]_net_1 , \sr_52_[9]_net_1 , \sr_52_[10]_net_1 , 
        \sr_52_[11]_net_1 , \sr_52_[12]_net_1 , \sr_51_[0]_net_1 , 
        \sr_51_[1]_net_1 , \sr_51_[2]_net_1 , \sr_51_[3]_net_1 , 
        \sr_51_[4]_net_1 , \sr_51_[5]_net_1 , \sr_51_[6]_net_1 , 
        \sr_51_[7]_net_1 , \sr_51_[8]_net_1 , \sr_51_[9]_net_1 , 
        \sr_51_[10]_net_1 , \sr_51_[11]_net_1 , \sr_51_[12]_net_1 , 
        \sr_50_[0]_net_1 , \sr_50_[1]_net_1 , \sr_50_[2]_net_1 , 
        \sr_50_[3]_net_1 , \sr_50_[4]_net_1 , \sr_50_[5]_net_1 , 
        \sr_50_[6]_net_1 , \sr_50_[7]_net_1 , \sr_50_[8]_net_1 , 
        \sr_50_[9]_net_1 , \sr_50_[10]_net_1 , \sr_50_[11]_net_1 , 
        \sr_50_[12]_net_1 , \sr_49_[0]_net_1 , \sr_49_[1]_net_1 , 
        \sr_49_[2]_net_1 , \sr_49_[3]_net_1 , \sr_49_[4]_net_1 , 
        \sr_49_[5]_net_1 , \sr_49_[6]_net_1 , \sr_49_[7]_net_1 , 
        \sr_49_[8]_net_1 , \sr_49_[9]_net_1 , \sr_49_[10]_net_1 , 
        \sr_49_[11]_net_1 , \sr_49_[12]_net_1 , \sr_48_[0]_net_1 , 
        \sr_48_[1]_net_1 , \sr_48_[2]_net_1 , \sr_48_[3]_net_1 , 
        \sr_48_[4]_net_1 , \sr_48_[5]_net_1 , \sr_48_[6]_net_1 , 
        \sr_48_[7]_net_1 , \sr_48_[8]_net_1 , \sr_48_[9]_net_1 , 
        \sr_48_[10]_net_1 , \sr_48_[11]_net_1 , \sr_48_[12]_net_1 , 
        \sr_47_[0]_net_1 , \sr_47_[1]_net_1 , \sr_47_[2]_net_1 , 
        \sr_47_[3]_net_1 , \sr_47_[4]_net_1 , \sr_47_[5]_net_1 , 
        \sr_47_[6]_net_1 , \sr_47_[7]_net_1 , \sr_47_[8]_net_1 , 
        \sr_47_[9]_net_1 , \sr_47_[10]_net_1 , \sr_47_[11]_net_1 , 
        \sr_47_[12]_net_1 , \sr_46_[0]_net_1 , \sr_46_[1]_net_1 , 
        \sr_46_[2]_net_1 , \sr_46_[3]_net_1 , \sr_46_[4]_net_1 , 
        \sr_46_[5]_net_1 , \sr_46_[6]_net_1 , \sr_46_[7]_net_1 , 
        \sr_46_[8]_net_1 , \sr_46_[9]_net_1 , \sr_46_[10]_net_1 , 
        \sr_46_[11]_net_1 , \sr_46_[12]_net_1 , \sr_45_[0]_net_1 , 
        \sr_45_[1]_net_1 , \sr_45_[2]_net_1 , \sr_45_[3]_net_1 , 
        \sr_45_[4]_net_1 , \sr_45_[5]_net_1 , \sr_45_[6]_net_1 , 
        \sr_45_[7]_net_1 , \sr_45_[8]_net_1 , \sr_45_[9]_net_1 , 
        \sr_45_[10]_net_1 , \sr_45_[11]_net_1 , \sr_45_[12]_net_1 , 
        \sr_44_[0]_net_1 , \sr_44_[1]_net_1 , \sr_44_[2]_net_1 , 
        \sr_44_[3]_net_1 , \sr_44_[4]_net_1 , \sr_44_[5]_net_1 , 
        \sr_44_[6]_net_1 , \sr_44_[7]_net_1 , \sr_44_[8]_net_1 , 
        \sr_44_[9]_net_1 , \sr_44_[10]_net_1 , \sr_44_[11]_net_1 , 
        \sr_44_[12]_net_1 , \sr_43_[0]_net_1 , \sr_43_[1]_net_1 , 
        \sr_43_[2]_net_1 , \sr_43_[3]_net_1 , \sr_43_[4]_net_1 , 
        \sr_43_[5]_net_1 , \sr_43_[6]_net_1 , \sr_43_[7]_net_1 , 
        \sr_43_[8]_net_1 , \sr_43_[9]_net_1 , \sr_43_[10]_net_1 , 
        \sr_43_[11]_net_1 , \sr_43_[12]_net_1 , \sr_42_[0]_net_1 , 
        \sr_42_[1]_net_1 , \sr_42_[2]_net_1 , \sr_42_[3]_net_1 , 
        \sr_42_[4]_net_1 , \sr_42_[5]_net_1 , \sr_42_[6]_net_1 , 
        \sr_42_[7]_net_1 , \sr_42_[8]_net_1 , \sr_42_[9]_net_1 , 
        \sr_42_[10]_net_1 , \sr_42_[11]_net_1 , \sr_42_[12]_net_1 , 
        \sr_41_[0]_net_1 , \sr_41_[1]_net_1 , \sr_41_[2]_net_1 , 
        \sr_41_[3]_net_1 , \sr_41_[4]_net_1 , \sr_41_[5]_net_1 , 
        \sr_41_[6]_net_1 , \sr_41_[7]_net_1 , \sr_41_[8]_net_1 , 
        \sr_41_[9]_net_1 , \sr_41_[10]_net_1 , \sr_41_[11]_net_1 , 
        \sr_41_[12]_net_1 , \sr_40_[0]_net_1 , \sr_40_[1]_net_1 , 
        \sr_40_[2]_net_1 , \sr_40_[3]_net_1 , \sr_40_[4]_net_1 , 
        \sr_40_[5]_net_1 , \sr_40_[6]_net_1 , \sr_40_[7]_net_1 , 
        \sr_40_[8]_net_1 , \sr_40_[9]_net_1 , \sr_40_[10]_net_1 , 
        \sr_40_[11]_net_1 , \sr_40_[12]_net_1 , \sr_62_[0]_net_1 , 
        \sr_62_[1]_net_1 , \sr_62_[2]_net_1 , \sr_62_[3]_net_1 , 
        \sr_62_[4]_net_1 , \sr_62_[5]_net_1 , \sr_62_[6]_net_1 , 
        \sr_62_[7]_net_1 , \sr_62_[8]_net_1 , \sr_62_[9]_net_1 , 
        \sr_62_[10]_net_1 , \sr_62_[11]_net_1 , \sr_62_[12]_net_1 , 
        \sr_61_[0]_net_1 , \sr_61_[1]_net_1 , \sr_61_[2]_net_1 , 
        \sr_61_[3]_net_1 , \sr_61_[4]_net_1 , \sr_61_[5]_net_1 , 
        \sr_61_[6]_net_1 , \sr_61_[7]_net_1 , \sr_61_[8]_net_1 , 
        \sr_61_[9]_net_1 , \sr_61_[10]_net_1 , \sr_61_[11]_net_1 , 
        \sr_61_[12]_net_1 , \sr_60_[0]_net_1 , \sr_60_[1]_net_1 , 
        \sr_60_[2]_net_1 , \sr_60_[3]_net_1 , \sr_60_[4]_net_1 , 
        \sr_60_[5]_net_1 , \sr_60_[6]_net_1 , \sr_60_[7]_net_1 , 
        \sr_60_[8]_net_1 , \sr_60_[9]_net_1 , \sr_60_[10]_net_1 , 
        \sr_60_[11]_net_1 , \sr_60_[12]_net_1 , \sr_59_[0]_net_1 , 
        \sr_59_[1]_net_1 , \sr_59_[2]_net_1 , \sr_59_[3]_net_1 , 
        \sr_59_[4]_net_1 , \sr_59_[5]_net_1 , \sr_59_[6]_net_1 , 
        \sr_59_[7]_net_1 , \sr_59_[8]_net_1 , \sr_59_[9]_net_1 , 
        \sr_59_[10]_net_1 , \sr_59_[11]_net_1 , \sr_59_[12]_net_1 , 
        \sr_58_[0]_net_1 , \sr_58_[1]_net_1 , \sr_58_[2]_net_1 , 
        \sr_58_[3]_net_1 , \sr_58_[4]_net_1 , \sr_58_[5]_net_1 , 
        \sr_58_[6]_net_1 , \sr_58_[7]_net_1 , \sr_58_[8]_net_1 , 
        \sr_58_[9]_net_1 , \sr_58_[10]_net_1 , \sr_58_[11]_net_1 , 
        \sr_58_[12]_net_1 , \sr_57_[0]_net_1 , \sr_57_[1]_net_1 , 
        \sr_57_[2]_net_1 , \sr_57_[3]_net_1 , \sr_57_[4]_net_1 , 
        \sr_57_[5]_net_1 , \sr_57_[6]_net_1 , \sr_57_[7]_net_1 , 
        \sr_57_[8]_net_1 , \sr_57_[9]_net_1 , \sr_57_[10]_net_1 , 
        \sr_57_[11]_net_1 , \sr_57_[12]_net_1 , \sr_56_[0]_net_1 , 
        \sr_56_[1]_net_1 , \sr_56_[2]_net_1 , \sr_56_[3]_net_1 , 
        \sr_56_[4]_net_1 , \sr_56_[5]_net_1 , \sr_56_[6]_net_1 , 
        \sr_56_[7]_net_1 , \sr_56_[8]_net_1 , \sr_56_[9]_net_1 , 
        \sr_56_[10]_net_1 , \sr_56_[11]_net_1 , \sr_56_[12]_net_1 , 
        \sr_55_[0]_net_1 , \sr_55_[1]_net_1 , \sr_55_[2]_net_1 , 
        \sr_55_[3]_net_1 , \sr_55_[4]_net_1 , \sr_55_[5]_net_1 , 
        \sr_55_[6]_net_1 , \sr_55_[7]_net_1 , \sr_55_[8]_net_1 , 
        \sr_55_[9]_net_1 , \sr_55_[10]_net_1 , \sr_55_[11]_net_1 , 
        \sr_55_[12]_net_1 , GND, VCC;
    
    DFN1E1C0 \sr_41_[5]  (.D(\sr_40_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[5]_net_1 ));
    DFN1E1C0 \sr_15_[3]  (.D(\sr_14_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[3]_net_1 ));
    DFN1E1C0 \sr_36_[5]  (.D(\sr_35_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[5]_net_1 ));
    DFN1E1C0 \sr_57_[5]  (.D(\sr_56_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[5]_net_1 ));
    DFN1E1C0 \sr_45_[11]  (.D(\sr_44_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[11]_net_1 ));
    DFN1E1C0 \sr_39_[6]  (.D(\sr_38_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[6]_net_1 ));
    DFN1E1C0 \sr_36_[4]  (.D(\sr_35_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[4]_net_1 ));
    DFN1E1C0 \sr_42_[4]  (.D(\sr_41_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[4]_net_1 ));
    DFN1E1C0 \sr_9_[3]  (.D(\sr_8_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[3]_net_1 ));
    DFN1E1C0 \sr_6_[4]  (.D(\sr_5_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[4]_net_1 ));
    DFN1E1C0 \sr_32_[3]  (.D(\sr_31_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[3]_net_1 ));
    DFN1E1C0 \sr_52_[6]  (.D(\sr_51_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[6]_net_1 ));
    DFN1E1C0 \sr_21_[9]  (.D(\sr_20_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[9]_net_1 ));
    DFN1E1C0 \sr_47_[12]  (.D(\sr_46_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[12]_net_1 ));
    DFN1E1C0 \sr_22_[4]  (.D(\sr_21_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[4]_net_1 ));
    DFN1E1C0 \sr_10_[1]  (.D(\sr_9_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[1]_net_1 ));
    DFN1E1C0 \sr_5_[4]  (.D(\sr_4_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[4]_net_1 ));
    DFN1E1C0 \sr_62_[6]  (.D(\sr_61_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[6]_net_1 ));
    DFN1E1C0 \sr_58_[2]  (.D(\sr_57_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[2]_net_1 ));
    DFN1E1C0 \sr_55_[0]  (.D(\sr_54_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[0]_net_1 ));
    DFN1E1C0 \sr_27_[3]  (.D(\sr_26_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[3]_net_1 ));
    DFN1E1C0 \sr_21_[1]  (.D(\sr_20_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[1]_net_1 ));
    DFN1E1C0 \sr_37_[9]  (.D(\sr_36_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[9]_net_1 ));
    DFN1E1C0 \sr_48_[10]  (.D(\sr_47_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[10]_net_1 ));
    DFN1E1C0 \sr_60_[5]  (.D(\sr_59_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[5]_net_1 ));
    DFN1E1C0 \sr_30_[5]  (.D(\sr_29_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[5]_net_1 ));
    DFN1E1C0 \sr_14_[4]  (.D(\sr_13_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[4]_net_1 ));
    DFN1E1C0 \sr_24_[8]  (.D(\sr_23_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[8]_net_1 ));
    DFN1E1C0 \sr_30_[4]  (.D(\sr_29_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[4]_net_1 ));
    DFN1E1C0 \sr_37_[6]  (.D(\sr_36_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[6]_net_1 ));
    DFN1E1C0 \sr_42_[6]  (.D(\sr_41_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[6]_net_1 ));
    DFN1E1C0 \sr_58_[4]  (.D(\sr_57_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[4]_net_1 ));
    DFN1E1C0 \sr_57_[10]  (.D(\sr_56_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[10]_net_1 ));
    DFN1E1C0 \sr_43_[7]  (.D(\sr_42_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[7]_net_1 ));
    DFN1E1C0 \sr_44_[2]  (.D(\sr_43_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[2]_net_1 ));
    DFN1E1C0 \sr_53_[7]  (.D(\sr_52_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[7]_net_1 ));
    DFN1E1C0 \sr_59_[1]  (.D(\sr_58_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[1]_net_1 ));
    DFN1E1C0 \sr_27_[10]  (.D(\sr_26_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[10]_net_1 ));
    DFN1E1C0 \sr_53_[8]  (.D(\sr_52_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[8]_net_1 ));
    DFN1E1C0 \sr_16_[4]  (.D(\sr_15_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[4]_net_1 ));
    DFN1E1C0 \sr_10_[11]  (.D(\sr_9_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[11]_net_1 ));
    DFN1E1C0 \sr_26_[8]  (.D(\sr_25_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[8]_net_1 ));
    DFN1E1C0 \sr_63_[7]  (.D(\sr_62_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[7]));
    DFN1E1C0 \sr_28_[7]  (.D(\sr_27_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[7]_net_1 ));
    DFN1E1C0 \sr_63_[8]  (.D(\sr_62_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[8]));
    DFN1E1C0 \sr_24_[0]  (.D(\sr_23_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[0]_net_1 ));
    DFN1E1C0 \sr_46_[2]  (.D(\sr_45_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[2]_net_1 ));
    DFN1E1C0 \sr_13_[5]  (.D(\sr_12_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[5]_net_1 ));
    DFN1E1C0 \sr_0_[2]  (.D(cur_error[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[2]));
    DFN1E1C0 \sr_0_[8]  (.D(cur_error[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[8]));
    DFN1E1C0 \sr_8_[3]  (.D(\sr_7_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[3]_net_1 ));
    DFN1E1C0 \sr_42_[11]  (.D(\sr_41_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[11]_net_1 ));
    DFN1E1C0 \sr_13_[3]  (.D(\sr_12_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[3]_net_1 ));
    DFN1E1C0 \sr_54_[10]  (.D(\sr_53_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[10]_net_1 ));
    DFN1E1C0 \sr_37_[11]  (.D(\sr_36_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[11]_net_1 ));
    DFN1E1C0 \sr_19_[7]  (.D(\sr_18_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[7]_net_1 ));
    DFN1E1C0 \sr_57_[1]  (.D(\sr_56_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[1]_net_1 ));
    DFN1E1C0 \sr_44_[11]  (.D(\sr_43_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[11]_net_1 ));
    DFN1E1C0 \sr_32_[10]  (.D(\sr_31_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[10]_net_1 ));
    DFN1E1C0 \sr_26_[0]  (.D(\sr_25_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[0]_net_1 ));
    DFN1E1C0 \sr_24_[10]  (.D(\sr_23_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[10]_net_1 ));
    DFN1E1C0 \sr_12_[1]  (.D(\sr_11_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[1]_net_1 ));
    DFN1E1C0 \sr_10_[4]  (.D(\sr_9_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[4]_net_1 ));
    DFN1E1C0 \sr_63_[0]  (.D(\sr_62_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[0]));
    DFN1E1C0 \sr_20_[8]  (.D(\sr_19_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[8]_net_1 ));
    DFN1E1C0 \sr_60_[12]  (.D(\sr_59_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[12]_net_1 ));
    DFN1E1C0 \sr_6_[10]  (.D(\sr_5_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[10]_net_1 ));
    DFN1E1C0 \sr_19_[6]  (.D(\sr_18_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[6]_net_1 ));
    DFN1E1C0 \sr_62_[5]  (.D(\sr_61_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[5]_net_1 ));
    DFN1E1C0 \sr_44_[8]  (.D(\sr_43_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[8]_net_1 ));
    DFN1E1C0 \sr_49_[5]  (.D(\sr_48_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[5]_net_1 ));
    DFN1E1C0 \sr_53_[0]  (.D(\sr_52_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[0]_net_1 ));
    DFN1E1C0 \sr_1_[2]  (.D(sr_new[2]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[2]));
    DFN1E1C0 \sr_40_[2]  (.D(\sr_39_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[2]_net_1 ));
    DFN1E1C0 \sr_32_[5]  (.D(\sr_31_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[5]_net_1 ));
    DFN1E1C0 \sr_1_[8]  (.D(sr_new[8]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[8]));
    DFN1E1C0 \sr_18_[12]  (.D(\sr_17_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[12]_net_1 ));
    DFN1E1C0 \sr_60_[10]  (.D(\sr_59_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[10]_net_1 ));
    DFN1E1C0 \sr_32_[4]  (.D(\sr_31_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[4]_net_1 ));
    DFN1E1C0 \sr_54_[3]  (.D(\sr_53_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[3]_net_1 ));
    DFN1E1C0 \sr_29_[9]  (.D(\sr_28_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[9]_net_1 ));
    DFN1E1C0 \sr_24_[2]  (.D(\sr_23_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[2]_net_1 ));
    DFN1E1C0 \sr_18_[9]  (.D(\sr_17_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[9]_net_1 ));
    DFN1E1C0 \sr_7_[9]  (.D(\sr_6_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[9]_net_1 ));
    DFN1E1C0 \sr_63_[10]  (.D(\sr_62_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[10]));
    DFN1E1C0 \sr_24_[5]  (.D(\sr_23_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[5]_net_1 ));
    DFN1E1C0 \sr_46_[8]  (.D(\sr_45_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[8]_net_1 ));
    DFN1E1C0 \sr_59_[11]  (.D(\sr_58_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[11]_net_1 ));
    DFN1E1C0 \sr_17_[7]  (.D(\sr_16_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[7]_net_1 ));
    DFN1E1C0 \sr_14_[8]  (.D(\sr_13_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[8]_net_1 ));
    DFN1E1C0 \sr_41_[3]  (.D(\sr_40_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[3]_net_1 ));
    DFN1E1C0 \sr_20_[0]  (.D(\sr_19_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[0]_net_1 ));
    DFN1E1C0 \sr_48_[0]  (.D(\sr_47_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[0]_net_1 ));
    DFN1E1C0 \sr_29_[1]  (.D(\sr_28_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[1]_net_1 ));
    DFN1E1C0 \sr_3_[10]  (.D(\sr_2_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[10]_net_1 ));
    DFN1E1C0 \sr_29_[11]  (.D(\sr_28_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[11]_net_1 ));
    DFN1E1C0 \sr_35_[1]  (.D(\sr_34_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[1]_net_1 ));
    DFN1E1C0 \sr_17_[6]  (.D(\sr_16_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[6]_net_1 ));
    DFN1E1C0 \sr_2_[3]  (.D(sr_prev[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[3]_net_1 ));
    DFN1E1C0 \sr_56_[3]  (.D(\sr_55_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[3]_net_1 ));
    DFN1E1C0 \sr_47_[5]  (.D(\sr_46_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[5]_net_1 ));
    DFN1E1C0 \sr_35_[2]  (.D(\sr_34_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[2]_net_1 ));
    DFN1E1C0 \sr_35_[12]  (.D(\sr_34_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[12]_net_1 ));
    DFN1E1C0 \sr_26_[2]  (.D(\sr_25_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[2]_net_1 ));
    DFN1E1C0 \sr_6_[2]  (.D(\sr_5_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[2]_net_1 ));
    DFN1E1C0 \sr_6_[8]  (.D(\sr_5_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[8]_net_1 ));
    DFN1E1C0 \sr_35_[7]  (.D(\sr_34_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[7]_net_1 ));
    DFN1E1C0 \sr_26_[5]  (.D(\sr_25_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[5]_net_1 ));
    DFN1E1C0 \sr_16_[8]  (.D(\sr_15_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[8]_net_1 ));
    DFN1E1C0 \sr_52_[12]  (.D(\sr_51_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[12]_net_1 ));
    DFN1E1C0 \sr_5_[2]  (.D(\sr_4_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[2]_net_1 ));
    DFN1E1C0 \sr_5_[8]  (.D(\sr_4_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[8]_net_1 ));
    DFN1E1C0 \sr_27_[9]  (.D(\sr_26_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[9]_net_1 ));
    DFN1E1C0 \sr_18_[11]  (.D(\sr_17_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[11]_net_1 ));
    DFN1E1C0 \sr_3_[9]  (.D(\sr_2_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[9]_net_1 ));
    DFN1E1C0 \sr_2_[11]  (.D(sr_prev[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[11]_net_1 ));
    DFN1E1C0 \sr_40_[8]  (.D(\sr_39_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[8]_net_1 ));
    DFN1E1C0 \sr_22_[12]  (.D(\sr_21_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[12]_net_1 ));
    DFN1E1C0 \sr_45_[9]  (.D(\sr_44_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[9]_net_1 ));
    DFN1E1C0 \sr_2_[12]  (.D(sr_prev[12]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[12]_net_1 ));
    DFN1E1C0 \sr_27_[1]  (.D(\sr_26_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[1]_net_1 ));
    DFN1E1C0 \sr_0__1[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_new_1_0));
    DFN1E1C0 \sr_9_[4]  (.D(\sr_8_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[4]_net_1 ));
    DFN1E1C0 \sr_12_[4]  (.D(\sr_11_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[4]_net_1 ));
    DFN1E1C0 \sr_56_[11]  (.D(\sr_55_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[11]_net_1 ));
    DFN1E1C0 \sr_22_[8]  (.D(\sr_21_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[8]_net_1 ));
    DFN1E1C0 \sr_14_[2]  (.D(\sr_13_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[2]_net_1 ));
    DFN1E1C0 \sr_46_[12]  (.D(\sr_45_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[12]_net_1 ));
    DFN1E1C0 \sr_50_[3]  (.D(\sr_49_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[3]_net_1 ));
    DFN1E1C0 \sr_20_[2]  (.D(\sr_19_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[2]_net_1 ));
    DFN1E1C0 \sr_44_[12]  (.D(\sr_43_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[12]_net_1 ));
    DFN1E1C0 \sr_26_[11]  (.D(\sr_25_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[11]_net_1 ));
    DFN1E1C0 \sr_14_[0]  (.D(\sr_13_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[0]_net_1 ));
    DFN1E1C0 \sr_34_[8]  (.D(\sr_33_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[8]_net_1 ));
    DFN1E1C0 \sr_20_[5]  (.D(\sr_19_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[5]_net_1 ));
    DFN1E1C0 \sr_10_[8]  (.D(\sr_9_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[8]_net_1 ));
    DFN1E1C0 \sr_42_[2]  (.D(\sr_41_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[2]_net_1 ));
    DFN1E1C0 \sr_55_[11]  (.D(\sr_54_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[11]_net_1 ));
    DFN1E1C0 \sr_51_[9]  (.D(\sr_50_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[9]_net_1 ));
    DFN1E1C0 \sr_54_[5]  (.D(\sr_53_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[5]_net_1 ));
    DFN1E1C0 \sr_25_[11]  (.D(\sr_24_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[11]_net_1 ));
    DFN1E1C0 \sr_21_[6]  (.D(\sr_20_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[6]_net_1 ));
    DFN1E1C0 \sr_57_[12]  (.D(\sr_56_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[12]_net_1 ));
    DFN1E1C0 \sr_16_[2]  (.D(\sr_15_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[2]_net_1 ));
    DFN1E1C0 \sr_35_[0]  (.D(\sr_34_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[0]_net_1 ));
    DFN1E1C0 \sr_16_[0]  (.D(\sr_15_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[0]_net_1 ));
    DFN1E1C0 \sr_36_[8]  (.D(\sr_35_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[8]_net_1 ));
    DFN1E1C0 \sr_27_[12]  (.D(\sr_26_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[12]_net_1 ));
    DFN1E1C0 \sr_22_[0]  (.D(\sr_21_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[0]_net_1 ));
    DFN1E1C0 \sr_0__0[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_new_0_0));
    DFN1E1C0 \sr_13_[11]  (.D(\sr_12_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[11]_net_1 ));
    DFN1E1C0 \sr_58_[10]  (.D(\sr_57_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[10]_net_1 ));
    DFN1E1C0 \sr_7_[12]  (.D(\sr_6_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[12]_net_1 ));
    DFN1E1C0 \sr_24_[3]  (.D(\sr_23_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[3]_net_1 ));
    DFN1E1C0 \sr_34_[9]  (.D(\sr_33_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[9]_net_1 ));
    DFN1E1C0 \sr_28_[10]  (.D(\sr_27_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[10]_net_1 ));
    DFN1E1C0 \sr_56_[5]  (.D(\sr_55_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[5]_net_1 ));
    DFN1E1C0 \sr_7_[10]  (.D(\sr_6_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[10]_net_1 ));
    DFN1E1C0 \sr_33_[1]  (.D(\sr_32_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[1]_net_1 ));
    DFN1E1C0 \sr_33_[2]  (.D(\sr_32_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[2]_net_1 ));
    DFN1E1C0 \sr_48_[7]  (.D(\sr_47_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[7]_net_1 ));
    DFN1E1C0 \sr_58_[7]  (.D(\sr_57_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[7]_net_1 ));
    DFN1E1C0 \sr_34_[6]  (.D(\sr_33_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[6]_net_1 ));
    DFN1E1C0 \sr_33_[7]  (.D(\sr_32_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[7]_net_1 ));
    DFN1E1C0 \sr_10_[2]  (.D(\sr_9_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[2]_net_1 ));
    DFN1E1C0 \sr_26_[3]  (.D(\sr_25_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[3]_net_1 ));
    DFN1E1C0 \sr_36_[9]  (.D(\sr_35_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[9]_net_1 ));
    DFN1E1C0 \sr_58_[8]  (.D(\sr_57_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[8]_net_1 ));
    DFN1E1C0 \sr_42_[8]  (.D(\sr_41_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[8]_net_1 ));
    DFN1E1C0 \sr_49_[3]  (.D(\sr_48_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[3]_net_1 ));
    DFN1E1C0 \sr_10_[0]  (.D(\sr_9_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[0]_net_1 ));
    DFN1E1C0 \sr_30_[8]  (.D(\sr_29_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[8]_net_1 ));
    DFN1E1C0 \sr_35_[10]  (.D(\sr_34_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[10]_net_1 ));
    DFN1E1C0 \sr_8_[4]  (.D(\sr_7_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[4]_net_1 ));
    DFN1E1C0 \sr_43_[12]  (.D(\sr_42_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[12]_net_1 ));
    DFN1E1C0 \sr_0_[9]  (.D(cur_error[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[9]));
    DFN1E1C0 \sr_43_[9]  (.D(\sr_42_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[9]_net_1 ));
    DFN1E1C0 \sr_50_[5]  (.D(\sr_49_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[5]_net_1 ));
    DFN1E1C0 \sr_52_[3]  (.D(\sr_51_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[3]_net_1 ));
    DFN1E1C0 \sr_22_[2]  (.D(\sr_21_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[2]_net_1 ));
    DFN1E1C0 \sr_18_[5]  (.D(\sr_17_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[5]_net_1 ));
    DFN1E1C0 \sr_7_[0]  (.D(\sr_6_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[0]_net_1 ));
    DFN1E1C0 \sr_36_[6]  (.D(\sr_35_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[6]_net_1 ));
    DFN1E1C0 \sr_60_[11]  (.D(\sr_59_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[11]_net_1 ));
    DFN1E1C0 \sr_45_[4]  (.D(\sr_44_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[4]_net_1 ));
    DFN1E1C0 \sr_22_[5]  (.D(\sr_21_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[5]_net_1 ));
    DFN1E1C0 \sr_35_[3]  (.D(\sr_34_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[3]_net_1 ));
    DFN1E1C0 \sr_7_[6]  (.D(\sr_6_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[6]_net_1 ));
    DFN1E1C0 \sr_12_[8]  (.D(\sr_11_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[8]_net_1 ));
    DFN1E1C0 \sr_55_[6]  (.D(\sr_54_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[6]_net_1 ));
    DFN1E1C0 \sr_52_[11]  (.D(\sr_51_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[11]_net_1 ));
    DFN1E1C0 \sr_18_[3]  (.D(\sr_17_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[3]_net_1 ));
    DFN1E1C0 \sr_36_[10]  (.D(\sr_35_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[10]_net_1 ));
    DFN1E1C0 \sr_25_[4]  (.D(\sr_24_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[4]_net_1 ));
    DFN1E1C0 \sr_22_[11]  (.D(\sr_21_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[11]_net_1 ));
    DFN1E1C0 \sr_20_[3]  (.D(\sr_19_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[3]_net_1 ));
    DFN1E1C0 \sr_30_[9]  (.D(\sr_29_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[9]_net_1 ));
    DFN1E1C0 \sr_47_[3]  (.D(\sr_46_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[3]_net_1 ));
    DFN1E1C0 \sr_54_[11]  (.D(\sr_53_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[11]_net_1 ));
    DFN1E1C0 \sr_4_[7]  (.D(\sr_3_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[7]_net_1 ));
    DFN1E1C0 \sr_31_[12]  (.D(\sr_30_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[12]_net_1 ));
    DFN1E1C0 \sr_54_[1]  (.D(\sr_53_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[1]_net_1 ));
    DFN1E1C0 \sr_24_[11]  (.D(\sr_23_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[11]_net_1 ));
    DFN1E1C0 \sr_1_[9]  (.D(sr_new[9]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[9]));
    DFN1E1C0 \sr_58_[0]  (.D(\sr_57_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[0]_net_1 ));
    DFN1E1C0 \sr_33_[0]  (.D(\sr_32_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[0]_net_1 ));
    DFN1E1C0 \sr_41_[1]  (.D(\sr_40_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[1]_net_1 ));
    DFN1E1C0 \sr_30_[6]  (.D(\sr_29_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[6]_net_1 ));
    DFN1E1C0 \sr_7_[1]  (.D(\sr_6_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[1]_net_1 ));
    DFN1E1C0 \sr_3_[0]  (.D(\sr_2_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[0]_net_1 ));
    DFN1E1C0 \sr_45_[6]  (.D(\sr_44_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[6]_net_1 ));
    DFN1E1C0 \sr_3_[6]  (.D(\sr_2_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[6]_net_1 ));
    DFN1E1C0 \sr_59_[9]  (.D(\sr_58_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[9]_net_1 ));
    DFN1E1C0 \sr_2_[4]  (.D(sr_prev[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[4]_net_1 ));
    DFN1E1C0 \sr_56_[1]  (.D(\sr_55_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[1]_net_1 ));
    DFN1E1C0 \sr_29_[6]  (.D(\sr_28_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[6]_net_1 ));
    DFN1E1C0 \sr_9_[2]  (.D(\sr_8_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[2]_net_1 ));
    DFN1E1C0 \sr_9_[8]  (.D(\sr_8_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[8]_net_1 ));
    DFN1E1C0 \sr_17_[11]  (.D(\sr_16_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[11]_net_1 ));
    DFN1E1C0 \sr_12_[2]  (.D(\sr_11_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[2]_net_1 ));
    DFN1E1C0 \sr_12_[10]  (.D(\sr_11_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[10]_net_1 ));
    DFN1E1C0 \sr_12_[0]  (.D(\sr_11_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[0]_net_1 ));
    DFN1E1C0 \sr_32_[8]  (.D(\sr_31_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[8]_net_1 ));
    DFN1E1C0 \sr_14_[7]  (.D(\sr_13_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[7]_net_1 ));
    DFN1E1C0 \sr_6_[9]  (.D(\sr_5_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[9]_net_1 ));
    DFN1E1C0 \sr_31_[10]  (.D(\sr_30_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[10]_net_1 ));
    DFN1E1C0 \sr_31_[11]  (.D(\sr_30_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[11]_net_1 ));
    DFN1E1C0 \sr_14_[6]  (.D(\sr_13_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[6]_net_1 ));
    DFN1E1C0 \sr_5_[10]  (.D(\sr_4_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[10]_net_1 ));
    DFN1E1C0 \sr_5_[9]  (.D(\sr_4_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[9]_net_1 ));
    DFN1E1C0 \sr_52_[5]  (.D(\sr_51_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[5]_net_1 ));
    DFN1E1C0 \sr_3_[1]  (.D(\sr_2_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[1]_net_1 ));
    DFN1E1C0 \sr_44_[5]  (.D(\sr_43_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[5]_net_1 ));
    DFN1E1C0 \sr_57_[9]  (.D(\sr_56_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[9]_net_1 ));
    DFN1E1C0 \sr_50_[1]  (.D(\sr_49_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[1]_net_1 ));
    DFN1E1C0 \sr_16_[7]  (.D(\sr_15_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[7]_net_1 ));
    DFN1E1C0 \sr_51_[2]  (.D(\sr_50_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[2]_net_1 ));
    DFN1E1C0 \sr_27_[6]  (.D(\sr_26_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[6]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1C0 \sr_43_[4]  (.D(\sr_42_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[4]_net_1 ));
    DFN1E1C0 \sr_24_[9]  (.D(\sr_23_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[9]_net_1 ));
    DFN1E1C0 \sr_22_[3]  (.D(\sr_21_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[3]_net_1 ));
    DFN1E1C0 \sr_33_[3]  (.D(\sr_32_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[3]_net_1 ));
    DFN1E1C0 \sr_32_[9]  (.D(\sr_31_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[9]_net_1 ));
    DFN1E1C0 \sr_15_[1]  (.D(\sr_14_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[1]_net_1 ));
    DFN1E1C0 \sr_53_[6]  (.D(\sr_52_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[6]_net_1 ));
    DFN1E1C0 \sr_60_[1]  (.D(\sr_59_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[1]_net_1 ));
    DFN1E1C0 \sr_16_[6]  (.D(\sr_15_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[6]_net_1 ));
    DFN1E1C0 \sr_61_[2]  (.D(\sr_60_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[2]_net_1 ));
    DFN1E1C0 \sr_23_[4]  (.D(\sr_22_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[4]_net_1 ));
    DFN1E1C0 \sr_46_[5]  (.D(\sr_45_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[5]_net_1 ));
    DFN1E1C0 \sr_24_[1]  (.D(\sr_23_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[1]_net_1 ));
    DFN1E1C0 \sr_63_[6]  (.D(\sr_62_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[6]));
    DFN1E1C0 \sr_49_[12]  (.D(\sr_48_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[12]_net_1 ));
    DFN1E1C0 \sr_56_[12]  (.D(\sr_55_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[12]_net_1 ));
    DFN1E1C0 \sr_54_[12]  (.D(\sr_53_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[12]_net_1 ));
    DFN1E1C0 \sr_35_[5]  (.D(\sr_34_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[5]_net_1 ));
    DFN1E1C0 \sr_15_[12]  (.D(\sr_14_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[12]_net_1 ));
    DFN1E1C0 \sr_32_[6]  (.D(\sr_31_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[6]_net_1 ));
    DFN1E1C0 \sr_26_[12]  (.D(\sr_25_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[12]_net_1 ));
    DFN1E1C0 \sr_35_[4]  (.D(\sr_34_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[4]_net_1 ));
    DFN1E1C0 \sr_26_[9]  (.D(\sr_25_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[9]_net_1 ));
    DFN1E1C0 \sr_24_[12]  (.D(\sr_23_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[12]_net_1 ));
    DFN1E1C0 \sr_51_[4]  (.D(\sr_50_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[4]_net_1 ));
    DFN1E1C0 \sr_10_[7]  (.D(\sr_9_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[7]_net_1 ));
    DFN1E1C0 \sr_8_[2]  (.D(\sr_7_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[2]_net_1 ));
    DFN1E1C0 \sr_40_[12]  (.D(\sr_39_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[12]_net_1 ));
    DFN1E1C0 \sr_8_[8]  (.D(\sr_7_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[8]_net_1 ));
    DFN1E1C0 \sr_26_[1]  (.D(\sr_25_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[1]_net_1 ));
    DFN1E1C0 \sr_61_[4]  (.D(\sr_60_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[4]_net_1 ));
    DFN1E1C0 \sr_0_[0]  (.D(cur_error[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[0]));
    DFN1E1C0 \sr_43_[6]  (.D(\sr_42_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[6]_net_1 ));
    DFN1E1C0 \sr_10_[6]  (.D(\sr_9_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[6]_net_1 ));
    DFN1E1C0 \sr_21_[7]  (.D(\sr_20_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[7]_net_1 ));
    DFN1E1C0 \sr_0_[6]  (.D(cur_error[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[6]));
    DFN1E1C0 \sr_40_[5]  (.D(\sr_39_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[5]_net_1 ));
    DFN1E1C0 \sr_40_[10]  (.D(\sr_39_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[10]_net_1 ));
    DFN1E1C0 \sr_43_[10]  (.D(\sr_42_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[10]_net_1 ));
    DFN1E1C0 \sr_38_[1]  (.D(\sr_37_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[1]_net_1 ));
    DFN1E1C0 \sr_49_[1]  (.D(\sr_48_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[1]_net_1 ));
    DFN1E1C0 \sr_63_[11]  (.D(\sr_62_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[11]));
    DFN1E1C0 \sr_20_[9]  (.D(\sr_19_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[9]_net_1 ));
    DFN1E1C0 \sr_38_[2]  (.D(\sr_37_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[2]_net_1 ));
    DFN1E1C0 \sr_38_[7]  (.D(\sr_37_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[7]_net_1 ));
    DFN1E1C0 \sr_52_[1]  (.D(\sr_51_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[1]_net_1 ));
    DFN1E1C0 \sr_20_[1]  (.D(\sr_19_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[1]_net_1 ));
    DFN1E1C0 \sr_1_[0]  (.D(sr_new[0]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[0]));
    DFN1E1C0 \sr_61_[9]  (.D(\sr_60_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[9]_net_1 ));
    DFN1E1C0 \sr_0_[1]  (.D(cur_error[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[1]));
    DFN1E1C0 \sr_15_[4]  (.D(\sr_14_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[4]_net_1 ));
    DFN1E1C0 \sr_1_[6]  (.D(sr_new[6]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[6]));
    DFN1E1C0 \sr_62_[1]  (.D(\sr_61_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[1]_net_1 ));
    DFN1E1C0 \sr_25_[8]  (.D(\sr_24_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[8]_net_1 ));
    DFN1E1C0 \sr_48_[9]  (.D(\sr_47_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[9]_net_1 ));
    DFN1E1C0 \sr_1_[11]  (.D(sr_new[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_prev[11]));
    DFN1E1C0 \sr_49_[10]  (.D(\sr_48_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[10]_net_1 ));
    DFN1E1C0 \sr_53_[12]  (.D(\sr_52_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[12]_net_1 ));
    DFN1E1C0 \sr_13_[1]  (.D(\sr_12_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[1]_net_1 ));
    DFN1E1C0 \sr_7_[5]  (.D(\sr_6_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[5]_net_1 ));
    DFN1E1C0 \sr_5_[12]  (.D(\sr_4_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[12]_net_1 ));
    DFN1E1C0 \sr_47_[1]  (.D(\sr_46_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[1]_net_1 ));
    DFN1E1C0 \sr_23_[12]  (.D(\sr_22_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[12]_net_1 ));
    DFN1E1C0 \sr_63_[5]  (.D(\sr_62_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[5]));
    DFN1E1C0 \sr_45_[2]  (.D(\sr_44_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[2]_net_1 ));
    DFN1E1C0 \sr_2_[2]  (.D(sr_prev[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[2]_net_1 ));
    DFN1E1C0 \sr_2_[8]  (.D(sr_prev[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[8]_net_1 ));
    DFN1E1C0 \sr_11_[9]  (.D(\sr_10_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[9]_net_1 ));
    DFN1E1C0 \sr_33_[5]  (.D(\sr_32_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[5]_net_1 ));
    DFN1E1C0 \sr_59_[2]  (.D(\sr_58_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[2]_net_1 ));
    DFN1E1C0 \sr_12_[7]  (.D(\sr_11_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[7]_net_1 ));
    DFN1E1C0 \sr_6_[0]  (.D(\sr_5_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[0]_net_1 ));
    DFN1E1C0 \sr_41_[0]  (.D(\sr_40_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[0]_net_1 ));
    DFN1E1C0 \sr_1_[1]  (.D(sr_new[1]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[1]));
    DFN1E1C0 \sr_33_[4]  (.D(\sr_32_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[4]_net_1 ));
    DFN1E1C0 \sr_9_[12]  (.D(\sr_8_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[12]_net_1 ));
    DFN1E1C0 \sr_25_[0]  (.D(\sr_24_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[0]_net_1 ));
    DFN1E1C0 \sr_6_[6]  (.D(\sr_5_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[6]_net_1 ));
    DFN1E1C0 \sr_15_[10]  (.D(\sr_14_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[10]_net_1 ));
    DFN1E1C0 \sr_12_[6]  (.D(\sr_11_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[6]_net_1 ));
    DFN1E1C0 \sr_61_[3]  (.D(\sr_60_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[3]_net_1 ));
    DFN1E1C0 \sr_5_[0]  (.D(\sr_4_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[0]_net_1 ));
    DFN1E1C0 \sr_44_[3]  (.D(\sr_43_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[3]_net_1 ));
    DFN1E1C0 \sr_38_[0]  (.D(\sr_37_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[0]_net_1 ));
    DFN1E1C0 \sr_42_[5]  (.D(\sr_41_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[5]_net_1 ));
    DFN1E1C0 \sr_5_[6]  (.D(\sr_4_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[6]_net_1 ));
    DFN1E1C0 \sr_3_[5]  (.D(\sr_2_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[5]_net_1 ));
    DFN1E1C0 \sr_4_[3]  (.D(\sr_3_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[3]_net_1 ));
    DFN1E1C0 \sr_9_[9]  (.D(\sr_8_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[9]_net_1 ));
    DFN1E1C0 \sr_37_[10]  (.D(\sr_36_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[10]_net_1 ));
    DFN1E1C0 \sr_22_[9]  (.D(\sr_21_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[9]_net_1 ));
    DFN1E1C0 \sr_59_[4]  (.D(\sr_58_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[4]_net_1 ));
    DFN1E1C0 \sr_16_[10]  (.D(\sr_15_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[10]_net_1 ));
    DFN1E1C0 \sr_57_[2]  (.D(\sr_56_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[2]_net_1 ));
    DFN1E1C0 \sr_46_[3]  (.D(\sr_45_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[3]_net_1 ));
    DFN1E1C0 \sr_6_[1]  (.D(\sr_5_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[1]_net_1 ));
    DFN1E1C0 \sr_45_[8]  (.D(\sr_44_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[8]_net_1 ));
    DFN1E1C0 \sr_22_[1]  (.D(\sr_21_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[1]_net_1 ));
    DFN1E1C0 \sr_29_[7]  (.D(\sr_28_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[7]_net_1 ));
    DFN1E1C0 \sr_11_[12]  (.D(\sr_10_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[12]_net_1 ));
    DFN1E1C0 \sr_5_[1]  (.D(\sr_4_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[1]_net_1 ));
    DFN1E1C0 \sr_4_[10]  (.D(\sr_3_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[10]_net_1 ));
    DFN1E1C0 \sr_55_[3]  (.D(\sr_54_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[3]_net_1 ));
    DFN1E1C0 \sr_25_[2]  (.D(\sr_24_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[2]_net_1 ));
    DFN1E1C0 \sr_13_[4]  (.D(\sr_12_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[4]_net_1 ));
    DFN1E1C0 \sr_62_[10]  (.D(\sr_61_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[10]_net_1 ));
    DFN1E1C0 \sr_23_[8]  (.D(\sr_22_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[8]_net_1 ));
    DFN1E1C0 \sr_25_[5]  (.D(\sr_24_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[5]_net_1 ));
    DFN1E1C0 \sr_15_[8]  (.D(\sr_14_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[8]_net_1 ));
    DFN1E1C0 \sr_34_[10]  (.D(\sr_33_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[10]_net_1 ));
    DFN1E1C0 \sr_57_[4]  (.D(\sr_56_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[4]_net_1 ));
    DFN1E1C0 \sr_40_[3]  (.D(\sr_39_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[3]_net_1 ));
    DFN1E1C0 \sr_48_[4]  (.D(\sr_47_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[4]_net_1 ));
    DFN1E1C0 \sr_38_[3]  (.D(\sr_37_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[3]_net_1 ));
    DFN1E1C0 \sr_43_[2]  (.D(\sr_42_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[2]_net_1 ));
    DFN1E1C0 \sr_58_[6]  (.D(\sr_57_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[6]_net_1 ));
    DFN1E1C0 \sr_54_[9]  (.D(\sr_53_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[9]_net_1 ));
    DFN1E1C0 \sr_28_[4]  (.D(\sr_27_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[4]_net_1 ));
    DFN1E1C0 \sr_27_[7]  (.D(\sr_26_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[7]_net_1 ));
    DFN1E1C0 \sr_24_[6]  (.D(\sr_23_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[6]_net_1 ));
    DFN1E1C0 \sr_40_[11]  (.D(\sr_39_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[11]_net_1 ));
    DFN1E1C0 \sr_11_[10]  (.D(\sr_10_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[10]_net_1 ));
    DFN1E1C0 \sr_23_[0]  (.D(\sr_22_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[0]_net_1 ));
    DFN1E1C0 \sr_11_[11]  (.D(\sr_10_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[11]_net_1 ));
    DFN1E1C0 \sr_59_[12]  (.D(\sr_58_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[12]_net_1 ));
    DFN1E1C0 \sr_8_[9]  (.D(\sr_7_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[9]_net_1 ));
    DFN1E1C0 \sr_1_[10]  (.D(sr_new[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_prev[10]));
    DFN1E1C0 \sr_41_[7]  (.D(\sr_40_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[7]_net_1 ));
    DFN1E1C0 \sr_29_[12]  (.D(\sr_28_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[12]_net_1 ));
    DFN1E1C0 \sr_19_[9]  (.D(\sr_18_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[9]_net_1 ));
    DFN1E1C0 \sr_56_[9]  (.D(\sr_55_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[9]_net_1 ));
    DFN1E1C0 \sr_51_[7]  (.D(\sr_50_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[7]_net_1 ));
    DFN1E1C0 \sr_39_[11]  (.D(\sr_38_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[11]_net_1 ));
    DFN1E1C0 \sr_26_[6]  (.D(\sr_25_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[6]_net_1 ));
    DFN1E1C0 \sr_51_[8]  (.D(\sr_50_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[8]_net_1 ));
    DFN1E1C0 \sr_50_[12]  (.D(\sr_49_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[12]_net_1 ));
    DFN1E1C0 \sr_49_[0]  (.D(\sr_48_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[0]_net_1 ));
    DFN1E1C0 \sr_0_[5]  (.D(cur_error[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[5]));
    DFN1E1C0 \sr_15_[2]  (.D(\sr_14_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[2]_net_1 ));
    DFN1E1C0 \sr_61_[7]  (.D(\sr_60_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[7]_net_1 ));
    DFN1E1C0 \sr_48_[6]  (.D(\sr_47_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[6]_net_1 ));
    DFN1E1C0 \sr_15_[0]  (.D(\sr_14_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[0]_net_1 ));
    DFN1E1C0 \sr_35_[8]  (.D(\sr_34_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[8]_net_1 ));
    DFN1E1C0 \sr_61_[8]  (.D(\sr_60_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[8]_net_1 ));
    DFN1E1C0 \sr_20_[12]  (.D(\sr_19_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[12]_net_1 ));
    DFN1E1C0 \sr_43_[8]  (.D(\sr_42_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[8]_net_1 ));
    DFN1E1C0 \sr_11_[5]  (.D(\sr_10_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[5]_net_1 ));
    DFN1E1C0 \sr_50_[10]  (.D(\sr_49_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[10]_net_1 ));
    DFN1E1C0 \sr_55_[5]  (.D(\sr_54_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[5]_net_1 ));
    DFN1E1C0 \sr_53_[10]  (.D(\sr_52_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[10]_net_1 ));
    DFN1E1C0 \sr_48_[12]  (.D(\sr_47_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[12]_net_1 ));
    DFN1E1C0 \sr_32_[12]  (.D(\sr_31_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[12]_net_1 ));
    DFN1E1C0 \sr_11_[3]  (.D(\sr_10_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[3]_net_1 ));
    DFN1E1C0 \sr_0_[11]  (.D(cur_error[11]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable), .Q(sr_new[11]));
    DFN1E1C0 \sr_20_[10]  (.D(\sr_19_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[10]_net_1 ));
    DFN1E1C0 \sr_50_[9]  (.D(\sr_49_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[9]_net_1 ));
    DFN1E1C0 \sr_17_[9]  (.D(\sr_16_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[9]_net_1 ));
    DFN1E1C0 \sr_23_[10]  (.D(\sr_22_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[10]_net_1 ));
    DFN1E1C0 \sr_20_[6]  (.D(\sr_19_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[6]_net_1 ));
    DFN1E1C0 \sr_53_[3]  (.D(\sr_52_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[3]_net_1 ));
    DFN1E1C0 \sr_23_[2]  (.D(\sr_22_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[2]_net_1 ));
    DFN1E1C0 \sr_1_[5]  (.D(sr_new[5]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[5]));
    DFN1E1C0 \sr_61_[0]  (.D(\sr_60_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[0]_net_1 ));
    DFN1E1C0 \sr_47_[0]  (.D(\sr_46_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[0]_net_1 ));
    DFN1E1C0 \sr_23_[5]  (.D(\sr_22_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[5]_net_1 ));
    DFN1E1C0 \sr_42_[3]  (.D(\sr_41_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[3]_net_1 ));
    DFN1E1C0 \sr_25_[3]  (.D(\sr_24_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[3]_net_1 ));
    DFN1E1C0 \sr_35_[9]  (.D(\sr_34_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[9]_net_1 ));
    DFN1E1C0 \sr_13_[8]  (.D(\sr_12_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[8]_net_1 ));
    DFN1E1C0 \sr_36_[11]  (.D(\sr_35_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[11]_net_1 ));
    DFN1E1C0 \sr_51_[0]  (.D(\sr_50_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[0]_net_1 ));
    DFN1E1C0 \sr_18_[1]  (.D(\sr_17_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[1]_net_1 ));
    DFN1E1C0 \sr_2_[9]  (.D(sr_prev[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[9]_net_1 ));
    DFN1E1C0 \sr_9_[0]  (.D(\sr_8_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[0]_net_1 ));
    DFN1E1C0 \sr_59_[10]  (.D(\sr_58_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[10]_net_1 ));
    DFN1E1C0 \sr_35_[11]  (.D(\sr_34_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[11]_net_1 ));
    DFN1E1C0 \sr_35_[6]  (.D(\sr_34_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[6]_net_1 ));
    DFN1E1C0 \sr_9_[6]  (.D(\sr_8_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[6]_net_1 ));
    DFN1E1C0 \sr_29_[10]  (.D(\sr_28_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[10]_net_1 ));
    DFN1E1C0 \sr_44_[1]  (.D(\sr_43_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[1]_net_1 ));
    DFN1E1C0 \sr_38_[5]  (.D(\sr_37_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[5]_net_1 ));
    DFN1E1C0 \sr_37_[12]  (.D(\sr_36_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[12]_net_1 ));
    DFN1E1C0 \sr_6_[5]  (.D(\sr_5_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[5]_net_1 ));
    DFN1E1C0 \sr_48_[11]  (.D(\sr_47_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[11]_net_1 ));
    DFN1E1C0 \sr_38_[4]  (.D(\sr_37_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[4]_net_1 ));
    DFN1E1C0 \sr_4_[4]  (.D(\sr_3_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[4]_net_1 ));
    DFN1E1C0 \sr_38_[10]  (.D(\sr_37_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[10]_net_1 ));
    DFN1E1C0 \sr_5_[5]  (.D(\sr_4_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[5]_net_1 ));
    DFN1E1C0 \sr_13_[2]  (.D(\sr_12_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[2]_net_1 ));
    DFN1E1C0 \sr_46_[1]  (.D(\sr_45_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[1]_net_1 ));
    DFN1E1C0 \sr_9_[1]  (.D(\sr_8_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[1]_net_1 ));
    DFN1E1C0 \sr_13_[0]  (.D(\sr_12_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[0]_net_1 ));
    DFN1E1C0 \sr_33_[8]  (.D(\sr_32_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[8]_net_1 ));
    DFN1E1C0 \sr_49_[7]  (.D(\sr_48_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[7]_net_1 ));
    DFN1E1C0 \sr_59_[7]  (.D(\sr_58_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[7]_net_1 ));
    DFN1E1C0 \sr_52_[9]  (.D(\sr_51_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[9]_net_1 ));
    DFN1E1C0 \sr_59_[8]  (.D(\sr_58_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[8]_net_1 ));
    DFN1E1C0 \sr_53_[5]  (.D(\sr_52_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[5]_net_1 ));
    DFN1E1C0 \sr_22_[6]  (.D(\sr_21_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[6]_net_1 ));
    DFN1E1C0 \sr_55_[1]  (.D(\sr_54_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[1]_net_1 ));
    DFN1E1C0 \sr_54_[2]  (.D(\sr_53_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[2]_net_1 ));
    DFN1E1C0 \sr_43_[11]  (.D(\sr_42_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[11]_net_1 ));
    DFN1E1C0 \sr_8_[0]  (.D(\sr_7_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[0]_net_1 ));
    DFN1E1C0 \sr_23_[3]  (.D(\sr_22_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[3]_net_1 ));
    DFN1E1C0 \sr_40_[1]  (.D(\sr_39_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[1]_net_1 ));
    DFN1E1C0 \sr_33_[9]  (.D(\sr_32_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[9]_net_1 ));
    DFN1E1C0 \sr_19_[5]  (.D(\sr_18_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[5]_net_1 ));
    DFN1E1C0 \sr_18_[4]  (.D(\sr_17_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[4]_net_1 ));
    DFN1E1C0 \sr_28_[8]  (.D(\sr_27_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[8]_net_1 ));
    DFN1E1C0 \sr_8_[6]  (.D(\sr_7_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[6]_net_1 ));
    DFN1E1C0 \sr_32_[11]  (.D(\sr_31_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[11]_net_1 ));
    DFN1E1C0 \sr_61_[12]  (.D(\sr_60_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[12]_net_1 ));
    DFN1E1C0 \sr_19_[3]  (.D(\sr_18_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[3]_net_1 ));
    DFN1E1C0 \sr_8_[11]  (.D(\sr_7_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[11]_net_1 ));
    DFN1E1C0 \sr_47_[7]  (.D(\sr_46_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[7]_net_1 ));
    DFN1E1C0 \sr_57_[7]  (.D(\sr_56_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[7]_net_1 ));
    DFN1E1C0 \sr_56_[2]  (.D(\sr_55_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[2]_net_1 ));
    DFN1E1C0 \sr_17_[10]  (.D(\sr_16_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[10]_net_1 ));
    DFN1E1C0 \sr_57_[8]  (.D(\sr_56_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[8]_net_1 ));
    DFN1E1C0 \sr_48_[2]  (.D(\sr_47_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[2]_net_1 ));
    DFN1E1C0 \sr_15_[7]  (.D(\sr_14_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[7]_net_1 ));
    DFN1E1C0 \sr_34_[11]  (.D(\sr_33_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[11]_net_1 ));
    DFN1E1C0 \sr_33_[6]  (.D(\sr_32_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[6]_net_1 ));
    DFN1E1C0 \sr_54_[4]  (.D(\sr_53_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[4]_net_1 ));
    DFN1E1C0 \sr_15_[6]  (.D(\sr_14_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[6]_net_1 ));
    DFN1E1C0 \sr_59_[0]  (.D(\sr_58_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[0]_net_1 ));
    DFN1E1C0 \sr_50_[11]  (.D(\sr_49_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[11]_net_1 ));
    DFN1E1C0 \sr_45_[5]  (.D(\sr_44_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[5]_net_1 ));
    DFN1E1C0 \sr_8_[1]  (.D(\sr_7_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[1]_net_1 ));
    DFN1E1C0 \sr_31_[1]  (.D(\sr_30_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[1]_net_1 ));
    DFN1E1C0 \sr_28_[0]  (.D(\sr_27_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[0]_net_1 ));
    DFN1E1C0 \sr_17_[5]  (.D(\sr_16_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[5]_net_1 ));
    DFN1E1C0 \sr_24_[7]  (.D(\sr_23_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[7]_net_1 ));
    DFN1E1C0 \sr_20_[11]  (.D(\sr_19_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[11]_net_1 ));
    DFN1E1C0 \sr_31_[2]  (.D(\sr_30_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[2]_net_1 ));
    DFN1E1C0 \sr_17_[3]  (.D(\sr_16_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[3]_net_1 ));
    DFN1E1C0 \sr_56_[4]  (.D(\sr_55_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[4]_net_1 ));
    DFN1E1C0 \sr_31_[7]  (.D(\sr_30_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[7]_net_1 ));
    DFN1E1C0 \sr_25_[9]  (.D(\sr_24_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[9]_net_1 ));
    DFN1E1C0 \sr_61_[10]  (.D(\sr_60_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[10]_net_1 ));
    DFN1E1C0 \sr_50_[2]  (.D(\sr_49_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[2]_net_1 ));
    DFN1E1C0 \sr_14_[10]  (.D(\sr_13_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[10]_net_1 ));
    DFN1E1C0 \sr_61_[11]  (.D(\sr_60_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[11]_net_1 ));
    DFN1E1C0 \sr_25_[1]  (.D(\sr_24_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[1]_net_1 ));
    DFN1E1C0 \sr_60_[2]  (.D(\sr_59_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[2]_net_1 ));
    DFN1E1C0 \sr_26_[7]  (.D(\sr_25_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[7]_net_1 ));
    DFN1E1C0 \sr_2_[0]  (.D(sr_prev[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[0]_net_1 ));
    DFN1E1C0 \sr_41_[9]  (.D(\sr_40_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[9]_net_1 ));
    DFN1E1C0 \sr_57_[0]  (.D(\sr_56_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[0]_net_1 ));
    DFN1E1C0 \sr_48_[8]  (.D(\sr_47_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[8]_net_1 ));
    DFN1E1C0 \sr_53_[1]  (.D(\sr_52_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[1]_net_1 ));
    DFN1E1C0 \sr_2_[6]  (.D(sr_prev[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[6]_net_1 ));
    DFN1E1C0 \sr_7_[7]  (.D(\sr_6_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[7]_net_1 ));
    DFN1E1C0 \sr_42_[1]  (.D(\sr_41_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[1]_net_1 ));
    DFN1E1C0 \sr_63_[1]  (.D(\sr_62_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[1]));
    DFN1E1C0 \sr_50_[4]  (.D(\sr_49_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[4]_net_1 ));
    DFN1E1C0 \sr_58_[12]  (.D(\sr_57_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[12]_net_1 ));
    DFN1E1C0 \sr_58_[3]  (.D(\sr_57_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[3]_net_1 ));
    DFN1E1C0 \sr_28_[2]  (.D(\sr_27_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[2]_net_1 ));
    DFN1E1C0 \sr_4_[2]  (.D(\sr_3_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[2]_net_1 ));
    DFN1E1C0 \sr_4_[8]  (.D(\sr_3_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[8]_net_1 ));
    DFN1E1C0 \sr_28_[5]  (.D(\sr_27_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[5]_net_1 ));
    DFN1E1C0 \sr_28_[12]  (.D(\sr_27_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[12]_net_1 ));
    DFN1E1C0 \sr_60_[4]  (.D(\sr_59_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[4]_net_1 ));
    DFN1E1C0 \sr_19_[11]  (.D(\sr_18_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[11]_net_1 ));
    DFN1E1C0 \sr_14_[9]  (.D(\sr_13_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[9]_net_1 ));
    DFN1E1C0 \sr_18_[8]  (.D(\sr_17_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[8]_net_1 ));
    DFN1E1C0 \sr_47_[11]  (.D(\sr_46_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[11]_net_1 ));
    DFN1E1C0 \sr_20_[7]  (.D(\sr_19_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[7]_net_1 ));
    DFN1E1C0 \sr_2_[1]  (.D(sr_prev[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[1]_net_1 ));
    DFN1E1C0 \sr_31_[0]  (.D(\sr_30_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[0]_net_1 ));
    DFN1E1C0 \sr_42_[10]  (.D(\sr_41_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[10]_net_1 ));
    DFN1E1C0 \sr_44_[0]  (.D(\sr_43_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[0]_net_1 ));
    DFN1E1C0 \sr_13_[7]  (.D(\sr_12_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[7]_net_1 ));
    DFN1E1C0 \sr_36_[12]  (.D(\sr_35_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[12]_net_1 ));
    DFN1E1C0 \sr_9_[5]  (.D(\sr_8_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[5]_net_1 ));
    DFN1E1C0 \sr_34_[12]  (.D(\sr_33_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[12]_net_1 ));
    DFN1E1C0 \sr_3_[7]  (.D(\sr_2_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[7]_net_1 ));
    DFN1E1C0 \sr_13_[6]  (.D(\sr_12_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[6]_net_1 ));
    DFN1E1C0 \sr_16_[9]  (.D(\sr_15_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[9]_net_1 ));
    DFN1E1C0 \sr_12_[12]  (.D(\sr_11_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[12]_net_1 ));
    DFN1E1C0 \sr_43_[5]  (.D(\sr_42_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[5]_net_1 ));
    DFN1E1C0 \sr_46_[0]  (.D(\sr_45_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[0]_net_1 ));
    DFN1E1C0 \sr_52_[2]  (.D(\sr_51_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[2]_net_1 ));
    DFN1E1C0 \sr_60_[9]  (.D(\sr_59_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[9]_net_1 ));
    DFN1E1C0 \sr_4_[12]  (.D(\sr_3_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[12]_net_1 ));
    DFN1E1C0 \sr_58_[11]  (.D(\sr_57_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[11]_net_1 ));
    DFN1E1C0 \sr_3_[12]  (.D(\sr_2_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[12]_net_1 ));
    DFN1E1C0 \sr_23_[9]  (.D(\sr_22_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[9]_net_1 ));
    DFN1E1C0 \sr_28_[11]  (.D(\sr_27_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[11]_net_1 ));
    DFN1E1C0 \sr_62_[2]  (.D(\sr_61_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[2]_net_1 ));
    DFN1E1C0 \sr_16_[11]  (.D(\sr_15_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[11]_net_1 ));
    DFN1E1C0 \sr_1_[12]  (.D(sr_new_0_0), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_prev[12]));
    DFN1E1C0 \sr_18_[2]  (.D(\sr_17_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[2]_net_1 ));
    DFN1E1C0 \sr_39_[1]  (.D(\sr_38_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[1]_net_1 ));
    DFN1E1C0 \sr_23_[1]  (.D(\sr_22_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[1]_net_1 ));
    DFN1E1C0 \sr_18_[0]  (.D(\sr_17_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[0]_net_1 ));
    DFN1E1C0 \sr_38_[8]  (.D(\sr_37_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[8]_net_1 ));
    DFN1E1C0 \sr_8_[10]  (.D(\sr_7_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[10]_net_1 ));
    DFN1E1C0 \sr_10_[9]  (.D(\sr_9_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[9]_net_1 ));
    DFN1E1C0 \sr_45_[12]  (.D(\sr_44_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[12]_net_1 ));
    DFN1E1C0 \sr_39_[2]  (.D(\sr_38_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[2]_net_1 ));
    DFN1E1C0 \sr_8_[12]  (.D(\sr_7_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[12]_net_1 ));
    DFN1E1C0 \sr_15_[11]  (.D(\sr_14_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[11]_net_1 ));
    DFN1E1C0 \sr_39_[7]  (.D(\sr_38_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[7]_net_1 ));
    DFN1E1C0 \sr_52_[4]  (.D(\sr_51_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[4]_net_1 ));
    DFN1E1C0 \sr_41_[4]  (.D(\sr_40_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[4]_net_1 ));
    DFN1E1C0 \sr_58_[5]  (.D(\sr_57_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[5]_net_1 ));
    DFN1E1C0 \sr_40_[0]  (.D(\sr_39_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[0]_net_1 ));
    DFN1E1C0 \sr_31_[3]  (.D(\sr_30_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[3]_net_1 ));
    DFN1E1C0 \sr_51_[6]  (.D(\sr_50_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[6]_net_1 ));
    DFN1E1C0 \sr_17_[12]  (.D(\sr_16_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[12]_net_1 ));
    DFN1E1C0 \sr_45_[3]  (.D(\sr_44_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[3]_net_1 ));
    DFN1E1C0 \sr_62_[4]  (.D(\sr_61_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[4]_net_1 ));
    DFN1E1C0 \sr_21_[4]  (.D(\sr_20_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[4]_net_1 ));
    DFN1E1C0 \sr_60_[3]  (.D(\sr_59_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[3]_net_1 ));
    DFN1E1C0 \sr_22_[7]  (.D(\sr_21_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[7]_net_1 ));
    DFN1E1C0 \sr_61_[6]  (.D(\sr_60_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[6]_net_1 ));
    DFN1E1C0 \sr_49_[9]  (.D(\sr_48_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[9]_net_1 ));
    DFN1E1C0 \sr_18_[10]  (.D(\sr_17_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[10]_net_1 ));
    DFN1E1C0 \sr_8_[5]  (.D(\sr_7_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[5]_net_1 ));
    DFN1E1C0 \sr_33_[12]  (.D(\sr_32_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[12]_net_1 ));
    DFN1E1C0 \sr_28_[3]  (.D(\sr_27_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[3]_net_1 ));
    DFN1E1C0 \sr_38_[9]  (.D(\sr_37_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[9]_net_1 ));
    DFN1E1C0 \sr_53_[11]  (.D(\sr_52_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[11]_net_1 ));
    DFN1E1C0 \sr_37_[1]  (.D(\sr_36_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[1]_net_1 ));
    DFN1E1C0 \sr_37_[2]  (.D(\sr_36_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[2]_net_1 ));
    DFN1E1C0 \sr_23_[11]  (.D(\sr_22_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[11]_net_1 ));
    DFN1E1C0 \sr_3_[11]  (.D(\sr_2_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[11]_net_1 ));
    DFN1E1C0 \sr_37_[7]  (.D(\sr_36_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[7]_net_1 ));
    DFN1E1C0 \sr_38_[6]  (.D(\sr_37_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[6]_net_1 ));
    DFN1E1C0 \sr_41_[6]  (.D(\sr_40_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[6]_net_1 ));
    DFN1E1C0 \sr_44_[7]  (.D(\sr_43_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[7]_net_1 ));
    DFN1E1C0 \sr_54_[7]  (.D(\sr_53_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[7]_net_1 ));
    DFN1E1C0 \sr_0_[7]  (.D(cur_error[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[7]));
    DFN1E1C0 \sr_9_[11]  (.D(\sr_8_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[11]_net_1 ));
    DFN1E1C0 \sr_62_[9]  (.D(\sr_61_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[9]_net_1 ));
    DFN1E1C0 \sr_54_[8]  (.D(\sr_53_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[8]_net_1 ));
    DFN1E1C0 \sr_39_[0]  (.D(\sr_38_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[0]_net_1 ));
    DFN1E1C0 \sr_47_[9]  (.D(\sr_46_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[9]_net_1 ));
    DFN1E1C0 \sr_6_[12]  (.D(\sr_5_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[12]_net_1 ));
    DFN1E1C0 \sr_7_[11]  (.D(\sr_6_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[11]_net_1 ));
    DFN1E1C0 \sr_46_[7]  (.D(\sr_45_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[7]_net_1 ));
    DFN1E1C0 \sr_14_[5]  (.D(\sr_13_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[5]_net_1 ));
    DFN1E1C0 \sr_56_[7]  (.D(\sr_55_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[7]_net_1 ));
    DFN1E1C0 \sr_12_[9]  (.D(\sr_11_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[9]_net_1 ));
    DFN1E1C0 \sr_12_[11]  (.D(\sr_11_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[11]_net_1 ));
    DFN1E1C0 \sr_55_[9]  (.D(\sr_54_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[9]_net_1 ));
    DFN1E1C0 \sr_56_[8]  (.D(\sr_55_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[8]_net_1 ));
    DFN1E1C0 \sr_25_[6]  (.D(\sr_24_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[6]_net_1 ));
    DFN1E1C0 \sr_14_[3]  (.D(\sr_13_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[3]_net_1 ));
    DFN1E1C0 \sr_42_[0]  (.D(\sr_41_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[0]_net_1 ));
    DFN1E1C0 \sr_1_[7]  (.D(sr_new[7]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[7]));
    DFN1E1C0 \sr_2_[5]  (.D(sr_prev[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[5]_net_1 ));
    DFN1E1C0 \sr_14_[11]  (.D(\sr_13_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[11]_net_1 ));
    DFN1E1C0 \sr_37_[0]  (.D(\sr_36_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[0]_net_1 ));
    DFN1E1C0 \sr_58_[1]  (.D(\sr_57_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[1]_net_1 ));
    DFN1E1C0 \sr_11_[1]  (.D(\sr_10_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[1]_net_1 ));
    DFN1E1C0 \sr_62_[3]  (.D(\sr_61_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[3]_net_1 ));
    DFN1E1C0 \sr_45_[10]  (.D(\sr_44_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[10]_net_1 ));
    DFN1E1C0 \sr_16_[5]  (.D(\sr_15_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[5]_net_1 ));
    DFN1E1C0 \sr_43_[3]  (.D(\sr_42_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[3]_net_1 ));
    DFN1E1C0 \sr_61_[5]  (.D(\sr_60_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[5]_net_1 ));
    DFN1E1C0 \sr_54_[0]  (.D(\sr_53_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[0]_net_1 ));
    DFN1E1C0 \sr_16_[3]  (.D(\sr_15_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[3]_net_1 ));
    DFN1E1C0 \sr_4_[9]  (.D(\sr_3_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[9]_net_1 ));
    DFN1E1C0 \sr_40_[7]  (.D(\sr_39_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[7]_net_1 ));
    DFN1E1C0 \sr_50_[7]  (.D(\sr_49_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[7]_net_1 ));
    DFN1E1C0 \sr_31_[5]  (.D(\sr_30_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[5]_net_1 ));
    DFN1E1C0 \sr_50_[8]  (.D(\sr_49_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[8]_net_1 ));
    DFN1E1C0 \sr_49_[4]  (.D(\sr_48_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[4]_net_1 ));
    DFN1E1C0 \sr_31_[4]  (.D(\sr_30_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[4]_net_1 ));
    DFN1E1C0 \sr_0_[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable), .Q(sr_new[12]));
    DFN1E1C0 \sr_39_[3]  (.D(\sr_38_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[3]_net_1 ));
    DFN1E1C0 \sr_6_[7]  (.D(\sr_5_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[7]_net_1 ));
    DFN1E1C0 \sr_60_[7]  (.D(\sr_59_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[7]_net_1 ));
    DFN1E1C0 \sr_59_[6]  (.D(\sr_58_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[6]_net_1 ));
    DFN1E1C0 \sr_7_[3]  (.D(\sr_6_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[3]_net_1 ));
    DFN1E1C0 \sr_46_[10]  (.D(\sr_45_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[10]_net_1 ));
    DFN1E1C0 \sr_60_[8]  (.D(\sr_59_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[8]_net_1 ));
    DFN1E1C0 \sr_29_[4]  (.D(\sr_28_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[4]_net_1 ));
    DFN1E1C0 \sr_57_[11]  (.D(\sr_56_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[11]_net_1 ));
    DFN1E1C0 \sr_56_[0]  (.D(\sr_55_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[0]_net_1 ));
    DFN1E1C0 \sr_5_[7]  (.D(\sr_4_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[7]_net_1 ));
    DFN1E1C0 \sr_18_[7]  (.D(\sr_17_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[7]_net_1 ));
    DFN1E1C0 \sr_10_[5]  (.D(\sr_9_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[5]_net_1 ));
    DFN1E1C0 \sr_41_[12]  (.D(\sr_40_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[12]_net_1 ));
    DFN1E1C0 \sr_52_[10]  (.D(\sr_51_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[10]_net_1 ));
    DFN1E1C0 \sr_27_[11]  (.D(\sr_26_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[11]_net_1 ));
    DFN1E1C0 \sr_39_[12]  (.D(\sr_38_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[12]_net_1 ));
    DFN1E1C0 \sr_18_[6]  (.D(\sr_17_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[6]_net_1 ));
    DFN1E1C0 \sr_22_[10]  (.D(\sr_21_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[10]_net_1 ));
    DFN1E1C0 \sr_10_[3]  (.D(\sr_9_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[3]_net_1 ));
    DFN1E1C0 \sr_48_[5]  (.D(\sr_47_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[5]_net_1 ));
    DFN1E1C0 \sr_60_[0]  (.D(\sr_59_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[0]_net_1 ));
    DFN1E1C0 \sr_47_[4]  (.D(\sr_46_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[4]_net_1 ));
    DFN1E1C0 \sr_30_[12]  (.D(\sr_29_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[12]_net_1 ));
    DFN1E1C0 \sr_37_[3]  (.D(\sr_36_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[3]_net_1 ));
    DFN1E1C0 \sr_57_[6]  (.D(\sr_56_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[6]_net_1 ));
    DFN1E1C0 \sr_49_[6]  (.D(\sr_48_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[6]_net_1 ));
    DFN1E1C0 \sr_3_[3]  (.D(\sr_2_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[3]_net_1 ));
    DFN1E1C0 \sr_28_[9]  (.D(\sr_27_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[9]_net_1 ));
    DFN1E1C0 \sr_27_[4]  (.D(\sr_26_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[4]_net_1 ));
    DFN1E1C0 \sr_62_[12]  (.D(\sr_61_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[12]_net_1 ));
    DFN1E1C0 \sr_50_[0]  (.D(\sr_49_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[0]_net_1 ));
    DFN1E1C0 \sr_53_[9]  (.D(\sr_52_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[9]_net_1 ));
    DFN1E1C0 \sr_23_[6]  (.D(\sr_22_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[6]_net_1 ));
    DFN1E1C0 \sr_28_[1]  (.D(\sr_27_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[1]_net_1 ));
    DFN1E1C0 \sr_11_[4]  (.D(\sr_10_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[4]_net_1 ));
    DFN1E1C0 \sr_30_[10]  (.D(\sr_29_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[10]_net_1 ));
    DFN1E1C0 \sr_21_[8]  (.D(\sr_20_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[8]_net_1 ));
    DFN1E1C0 \sr_16_[12]  (.D(\sr_15_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[12]_net_1 ));
    DFN1E1C0 \sr_41_[10]  (.D(\sr_40_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[10]_net_1 ));
    DFN1E1C0 \sr_45_[1]  (.D(\sr_44_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[1]_net_1 ));
    DFN1E1C0 \sr_33_[10]  (.D(\sr_32_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[10]_net_1 ));
    DFN1E1C0 \sr_14_[12]  (.D(\sr_13_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[12]_net_1 ));
    DFN1E1C0 \sr_41_[11]  (.D(\sr_40_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[11]_net_1 ));
    DFN1E1C0 \sr_55_[12]  (.D(\sr_54_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[12]_net_1 ));
    DFN1E1C0 \sr_42_[7]  (.D(\sr_41_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[7]_net_1 ));
    DFN1E1C0 \sr_52_[7]  (.D(\sr_51_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[7]_net_1 ));
    DFN1E1C0 \sr_41_[2]  (.D(\sr_40_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[2]_net_1 ));
    DFN1E1C0 \sr_52_[8]  (.D(\sr_51_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[8]_net_1 ));
    DFN1E1C0 \sr_25_[12]  (.D(\sr_24_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[12]_net_1 ));
    DFN1E1C0 \sr_47_[6]  (.D(\sr_46_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[6]_net_1 ));
    DFN1E1C0 \sr_62_[7]  (.D(\sr_61_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[7]_net_1 ));
    DFN1E1C0 \sr_62_[8]  (.D(\sr_61_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[8]_net_1 ));
    DFN1E1C0 \sr_19_[1]  (.D(\sr_18_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[1]_net_1 ));
    DFN1E1C0 \sr_21_[0]  (.D(\sr_20_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[0]_net_1 ));
    DFN1E1C0 \sr_39_[10]  (.D(\sr_38_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[10]_net_1 ));
    DFN1E1C0 \sr_12_[5]  (.D(\sr_11_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[5]_net_1 ));
    DFN1E1C0 \sr_0_[10]  (.D(cur_error[10]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable), .Q(sr_new[10]));
    DFN1E1C0 \sr_12_[3]  (.D(\sr_11_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[3]_net_1 ));
    DFN1E1C0 \sr_34_[1]  (.D(\sr_33_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[1]_net_1 ));
    DFN1E1C0 \sr_39_[5]  (.D(\sr_38_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[5]_net_1 ));
    DFN1E1C0 \sr_5_[11]  (.D(\sr_4_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[11]_net_1 ));
    DFN1E1C0 \sr_34_[2]  (.D(\sr_33_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[2]_net_1 ));
    DFN1E1C0 \sr_39_[4]  (.D(\sr_38_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[4]_net_1 ));
    DFN1E1C0 \sr_55_[2]  (.D(\sr_54_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[2]_net_1 ));
    DFN1E1C0 \sr_62_[0]  (.D(\sr_61_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[0]_net_1 ));
    DFN1E1C0 \sr_34_[7]  (.D(\sr_33_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[7]_net_1 ));
    DFN1E1C0 \sr_41_[8]  (.D(\sr_40_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[8]_net_1 ));
    DFN1E1C0 \sr_52_[0]  (.D(\sr_51_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[0]_net_1 ));
    DFN1E1C0 \sr_17_[1]  (.D(\sr_16_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[1]_net_1 ));
    DFN1E1C0 \sr_4_[0]  (.D(\sr_3_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[0]_net_1 ));
    DFN1E1C0 \sr_36_[1]  (.D(\sr_35_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[1]_net_1 ));
    DFN1E1C0 \sr_13_[12]  (.D(\sr_12_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[12]_net_1 ));
    DFN1E1C0 \sr_4_[6]  (.D(\sr_3_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[6]_net_1 ));
    DFN1E1C0 \sr_44_[9]  (.D(\sr_43_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[9]_net_1 ));
    DFN1E1C0 \sr_0_[3]  (.D(cur_error[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[3]));
    DFN1E1C0 \sr_36_[2]  (.D(\sr_35_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[2]_net_1 ));
    DFN1E1C0 \sr_51_[3]  (.D(\sr_50_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[3]_net_1 ));
    DFN1E1C0 \sr_36_[7]  (.D(\sr_35_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[7]_net_1 ));
    DFN1E1C0 \sr_21_[2]  (.D(\sr_20_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[2]_net_1 ));
    DFN1E1C0 \sr_37_[5]  (.D(\sr_36_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[5]_net_1 ));
    DFN1E1C0 \sr_55_[4]  (.D(\sr_54_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[4]_net_1 ));
    DFN1E1C0 \sr_21_[5]  (.D(\sr_20_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[5]_net_1 ));
    DFN1E1C0 \sr_43_[1]  (.D(\sr_42_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[1]_net_1 ));
    DFN1E1C0 \sr_11_[8]  (.D(\sr_10_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[8]_net_1 ));
    DFN1E1C0 \sr_37_[4]  (.D(\sr_36_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[4]_net_1 ));
    DFN1E1C0 \sr_62_[11]  (.D(\sr_61_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[11]_net_1 ));
    DFN1E1C0 \sr_46_[9]  (.D(\sr_45_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[9]_net_1 ));
    DFN1E1C0 \sr_25_[7]  (.D(\sr_24_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[7]_net_1 ));
    DFN1E1C0 \sr_48_[3]  (.D(\sr_47_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[3]_net_1 ));
    DFN1E1C0 \sr_30_[1]  (.D(\sr_29_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[1]_net_1 ));
    DFN1E1C0 \sr_4_[1]  (.D(\sr_3_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[1]_net_1 ));
    DFN1E1C0 \sr_55_[10]  (.D(\sr_54_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[10]_net_1 ));
    DFN1E1C0 \sr_19_[4]  (.D(\sr_18_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[4]_net_1 ));
    DFN1E1C0 \sr_9_[7]  (.D(\sr_8_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[7]_net_1 ));
    DFN1E1C0 \sr_7_[4]  (.D(\sr_6_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[4]_net_1 ));
    DFN1E1C0 \sr_29_[8]  (.D(\sr_28_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[8]_net_1 ));
    DFN1E1C0 \sr_1_[3]  (.D(sr_new[3]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[3]));
    DFN1E1C0 \sr_34_[0]  (.D(\sr_33_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[0]_net_1 ));
    DFN1E1C0 \sr_30_[2]  (.D(\sr_29_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[2]_net_1 ));
    DFN1E1C0 \sr_25_[10]  (.D(\sr_24_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[10]_net_1 ));
    DFN1E1C0 \sr_30_[7]  (.D(\sr_29_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[7]_net_1 ));
    DFN1E1C0 \sr_49_[2]  (.D(\sr_48_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[2]_net_1 ));
    DFN1E1C0 \sr_56_[10]  (.D(\sr_55_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[10]_net_1 ));
    DFN1E1C0 \sr_40_[9]  (.D(\sr_39_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[9]_net_1 ));
    DFN1E1C0 \sr_36_[0]  (.D(\sr_35_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[0]_net_1 ));
    DFN1E1C0 \sr_11_[2]  (.D(\sr_10_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[2]_net_1 ));
    DFN1E1C0 \sr_30_[11]  (.D(\sr_29_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[11]_net_1 ));
    DFN1E1C0 \sr_53_[2]  (.D(\sr_52_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[2]_net_1 ));
    DFN1E1C0 \sr_26_[10]  (.D(\sr_25_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[10]_net_1 ));
    DFN1E1C0 \sr_11_[0]  (.D(\sr_10_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[0]_net_1 ));
    DFN1E1C0 \sr_31_[8]  (.D(\sr_30_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[8]_net_1 ));
    DFN1E1C0 \sr_29_[0]  (.D(\sr_28_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[0]_net_1 ));
    DFN1E1C0 \sr_17_[4]  (.D(\sr_16_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[4]_net_1 ));
    DFN1E1C0 \sr_6_[3]  (.D(\sr_5_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[3]_net_1 ));
    DFN1E1C0 \sr_51_[12]  (.D(\sr_50_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[12]_net_1 ));
    DFN1E1C0 \sr_27_[8]  (.D(\sr_26_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[8]_net_1 ));
    DFN1E1C0 \sr_3_[4]  (.D(\sr_2_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[4]_net_1 ));
    DFN1E1C0 \sr_63_[2]  (.D(\sr_62_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[2]));
    DFN1E1C0 \sr_21_[12]  (.D(\sr_20_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[12]_net_1 ));
    DFN1E1C0 \sr_5_[3]  (.D(\sr_4_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[3]_net_1 ));
    DFN1E1C0 \sr_15_[9]  (.D(\sr_14_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[9]_net_1 ));
    DFN1E1C0 \sr_51_[5]  (.D(\sr_50_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[5]_net_1 ));
    DFN1E1C0 \sr_47_[2]  (.D(\sr_46_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[2]_net_1 ));
    DFN1E1C0 \sr_47_[10]  (.D(\sr_46_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[10]_net_1 ));
    DFN1E1C0 \sr_45_[0]  (.D(\sr_44_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[0]_net_1 ));
    DFN1E1C0 \sr_58_[9]  (.D(\sr_57_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[9]_net_1 ));
    DFN1E1C0 \sr_30_[0]  (.D(\sr_29_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[0]_net_1 ));
    DFN1E1C0 \sr_44_[4]  (.D(\sr_43_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[4]_net_1 ));
    DFN1E1C0 \sr_53_[4]  (.D(\sr_52_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[4]_net_1 ));
    DFN1E1C0 \sr_34_[3]  (.D(\sr_33_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[3]_net_1 ));
    DFN1E1C0 \sr_54_[6]  (.D(\sr_53_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[6]_net_1 ));
    DFN1E1C0 \sr_49_[8]  (.D(\sr_48_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[8]_net_1 ));
    DFN1E1C0 \sr_28_[6]  (.D(\sr_27_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[6]_net_1 ));
    DFN1E1C0 \sr_21_[3]  (.D(\sr_20_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[3]_net_1 ));
    DFN1E1C0 \sr_31_[9]  (.D(\sr_30_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[9]_net_1 ));
    DFN1E1C0 \sr_8_[7]  (.D(\sr_7_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[7]_net_1 ));
    DFN1E1C0 \sr_27_[0]  (.D(\sr_26_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[0]_net_1 ));
    DFN1E1C0 \sr_24_[4]  (.D(\sr_23_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[4]_net_1 ));
    DFN1E1C0 \sr_63_[4]  (.D(\sr_62_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[4]));
    DFN1E1C0 \sr_32_[1]  (.D(\sr_31_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[1]_net_1 ));
    DFN1E1C0 \sr_19_[12]  (.D(\sr_18_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[12]_net_1 ));
    DFN1E1C0 \sr_23_[7]  (.D(\sr_22_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[7]_net_1 ));
    DFN1E1C0 \sr_51_[10]  (.D(\sr_50_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[10]_net_1 ));
    DFN1E1C0 \sr_32_[2]  (.D(\sr_31_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[2]_net_1 ));
    DFN1E1C0 \sr_38_[12]  (.D(\sr_37_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[12]_net_1 ));
    DFN1E1C0 \sr_59_[3]  (.D(\sr_58_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[3]_net_1 ));
    DFN1E1C0 \sr_51_[11]  (.D(\sr_50_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[11]_net_1 ));
    DFN1E1C0 \sr_29_[2]  (.D(\sr_28_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[2]_net_1 ));
    DFN1E1C0 \sr_32_[7]  (.D(\sr_31_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[7]_net_1 ));
    DFN1E1C0 \sr_21_[10]  (.D(\sr_20_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[10]_net_1 ));
    DFN1E1C0 \sr_46_[4]  (.D(\sr_45_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[4]_net_1 ));
    DFN1E1C0 \sr_31_[6]  (.D(\sr_30_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[6]_net_1 ));
    DFN1E1C0 \sr_36_[3]  (.D(\sr_35_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[3]_net_1 ));
    DFN1E1C0 \sr_29_[5]  (.D(\sr_28_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[5]_net_1 ));
    DFN1E1C0 \sr_56_[6]  (.D(\sr_55_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[6]_net_1 ));
    DFN1E1C0 \sr_21_[11]  (.D(\sr_20_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[11]_net_1 ));
    DFN1E1C0 \sr_19_[8]  (.D(\sr_18_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[8]_net_1 ));
    DFN1E1C0 \sr_44_[10]  (.D(\sr_43_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[10]_net_1 ));
    DFN1E1C0 \sr_10_[12]  (.D(\sr_9_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[12]_net_1 ));
    DFN1E1C0 \sr_26_[4]  (.D(\sr_25_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[4]_net_1 ));
    DFN1E1C0 \sr_47_[8]  (.D(\sr_46_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[8]_net_1 ));
    DFN1E1C0 \sr_44_[6]  (.D(\sr_43_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[6]_net_1 ));
    DFN1E1C0 \sr_42_[9]  (.D(\sr_41_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[9]_net_1 ));
    DFN1E1C0 \sr_63_[9]  (.D(\sr_62_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[9]));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \sr_10_[10]  (.D(\sr_9_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[10]_net_1 ));
    DFN1E1C0 \sr_2_[10]  (.D(sr_prev[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[10]_net_1 ));
    DFN1E1C0 \sr_13_[10]  (.D(\sr_12_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[10]_net_1 ));
    DFN1E1C0 \sr_57_[3]  (.D(\sr_56_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[3]_net_1 ));
    DFN1E1C0 \sr_27_[2]  (.D(\sr_26_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[2]_net_1 ));
    DFN1E1C0 \sr_40_[4]  (.D(\sr_39_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[4]_net_1 ));
    DFN1E1C0 \sr_30_[3]  (.D(\sr_29_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[3]_net_1 ));
    DFN1E1C0 \sr_50_[6]  (.D(\sr_49_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[6]_net_1 ));
    DFN1E1C0 \sr_27_[5]  (.D(\sr_26_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[5]_net_1 ));
    DFN1E1C0 \sr_46_[6]  (.D(\sr_45_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[6]_net_1 ));
    DFN1E1C0 \sr_38_[11]  (.D(\sr_37_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[11]_net_1 ));
    DFN1E1C0 \sr_17_[8]  (.D(\sr_16_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[8]_net_1 ));
    DFN1E1C0 \sr_20_[4]  (.D(\sr_19_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[4]_net_1 ));
    DFN1E1C0 \sr_0_[4]  (.D(cur_error[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[4]));
    DFN1E1C0 \sr_49_[11]  (.D(\sr_48_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[11]_net_1 ));
    DFN1E1C0 \sr_13_[9]  (.D(\sr_12_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[9]_net_1 ));
    DFN1E1C0 \sr_60_[6]  (.D(\sr_59_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[6]_net_1 ));
    DFN1E1C0 \sr_2_[7]  (.D(sr_prev[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[7]_net_1 ));
    DFN1E1C0 \sr_51_[1]  (.D(\sr_50_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[1]_net_1 ));
    DFN1E1C0 \sr_32_[0]  (.D(\sr_31_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[0]_net_1 ));
    DFN1E1C0 \sr_7_[2]  (.D(\sr_6_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[2]_net_1 ));
    DFN1E1C0 \sr_4_[11]  (.D(\sr_3_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[11]_net_1 ));
    DFN1E1C0 \sr_19_[2]  (.D(\sr_18_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[2]_net_1 ));
    DFN1E1C0 \sr_7_[8]  (.D(\sr_6_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[8]_net_1 ));
    DFN1E1C0 \sr_4_[5]  (.D(\sr_3_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[5]_net_1 ));
    DFN1E1C0 \sr_43_[0]  (.D(\sr_42_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[0]_net_1 ));
    DFN1E1C0 \sr_19_[0]  (.D(\sr_18_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[0]_net_1 ));
    DFN1E1C0 \sr_9_[10]  (.D(\sr_8_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[10]_net_1 ));
    DFN1E1C0 \sr_39_[8]  (.D(\sr_38_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[8]_net_1 ));
    DFN1E1C0 \sr_61_[1]  (.D(\sr_60_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[1]_net_1 ));
    DFN1E1C0 \sr_19_[10]  (.D(\sr_18_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[10]_net_1 ));
    DFN1E1C0 \sr_14_[1]  (.D(\sr_13_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[1]_net_1 ));
    DFN1E1C0 \sr_63_[3]  (.D(\sr_62_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[3]));
    DFN1E1C0 \sr_45_[7]  (.D(\sr_44_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[7]_net_1 ));
    DFN1E1C0 \sr_59_[5]  (.D(\sr_58_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[5]_net_1 ));
    DFN1E1C0 \sr_55_[7]  (.D(\sr_54_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[7]_net_1 ));
    DFN1E1C0 \sr_63_[12]  (.D(\sr_62_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[12]));
    DFN1E1C0 \sr_48_[1]  (.D(\sr_47_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[1]_net_1 ));
    DFN1E1C0 \sr_42_[12]  (.D(\sr_41_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[12]_net_1 ));
    DFN1E1C0 \sr_40_[6]  (.D(\sr_39_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[6]_net_1 ));
    DFN1E1C0 \sr_55_[8]  (.D(\sr_54_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[8]_net_1 ));
    DFN1E1C0 \sr_1_[4]  (.D(sr_new[4]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[4]));
    DFN1E1C0 \sr_34_[5]  (.D(\sr_33_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[5]_net_1 ));
    DFN1E1C0 \sr_6_[11]  (.D(\sr_5_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[11]_net_1 ));
    DFN1E1C0 \sr_11_[7]  (.D(\sr_10_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[7]_net_1 ));
    DFN1E1C0 \sr_34_[4]  (.D(\sr_33_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[4]_net_1 ));
    DFN1E1C0 \sr_16_[1]  (.D(\sr_15_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[1]_net_1 ));
    DFN1E1C0 \sr_29_[3]  (.D(\sr_28_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[3]_net_1 ));
    DFN1E1C0 \sr_17_[2]  (.D(\sr_16_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[2]_net_1 ));
    DFN1E1C0 \sr_39_[9]  (.D(\sr_38_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[9]_net_1 ));
    DFN1E1C0 \sr_3_[2]  (.D(\sr_2_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[2]_net_1 ));
    DFN1E1C0 \sr_46_[11]  (.D(\sr_45_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[11]_net_1 ));
    DFN1E1C0 \sr_3_[8]  (.D(\sr_2_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[8]_net_1 ));
    DFN1E1C0 \sr_33_[11]  (.D(\sr_32_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[11]_net_1 ));
    DFN1E1C0 \sr_17_[0]  (.D(\sr_16_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[0]_net_1 ));
    DFN1E1C0 \sr_37_[8]  (.D(\sr_36_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[8]_net_1 ));
    DFN1E1C0 \sr_15_[5]  (.D(\sr_14_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[5]_net_1 ));
    DFN1E1C0 \sr_11_[6]  (.D(\sr_10_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[6]_net_1 ));
    
endmodule


module controller_Z1_4_2(
       state_0_0,
       state_0_d0,
       pwm_chg,
       sig_prev,
       sig_old_i_0,
       avg_done,
       N_46_1,
       vd_rdy,
       sum_rdy,
       deriv_enable,
       calc_avg,
       calc_int,
       pwm_enable,
       sum_enable,
       calc_error,
       avg_enable,
       int_enable,
       pwm_chg_0,
       avg_enable_0,
       n_rst_c,
       clk_c,
       avg_enable_1
    );
input  state_0_0;
input  state_0_d0;
output pwm_chg;
input  sig_prev;
input  sig_old_i_0;
input  avg_done;
input  N_46_1;
input  vd_rdy;
input  sum_rdy;
output deriv_enable;
output calc_avg;
output calc_int;
output pwm_enable;
output sum_enable;
output calc_error;
output avg_enable;
output int_enable;
output pwm_chg_0;
output avg_enable_0;
input  n_rst_c;
input  clk_c;
output avg_enable_1;

    wire \state_RNI808O1[0]_net_1 , N_12, \state_0[5] , N_94, 
        \count[13]_net_1 , count_c12, count_31_0, count_n14, 
        count_n14_tz, N_62, \count[14]_net_1 , count_n13, count_n11, 
        count_c10, \count[11]_net_1 , count_n12, count_c11, 
        \count[12]_net_1 , count_n15, \count[15]_net_1 , count_c7, 
        count_c6, \count[7]_net_1 , count_c5, \count[6]_net_1 , 
        count_c4, \count[5]_net_1 , count_c3, \count[4]_net_1 , 
        count_c2, \count[3]_net_1 , count_c1, \count[2]_net_1 , 
        \count[0]_net_1 , \count[1]_net_1 , count_c8, \count[8]_net_1 , 
        count_c9, \count[9]_net_1 , \count[10]_net_1 , 
        \state_ns_0_a2_9[0] , \state[10]_net_1 , N_33, 
        \state_ns_0_a2_8[0] , \state_ns_0_a2_6[0] , 
        \state_ns_0_a2_5[0] , \state_ns_0_a2_2[0] , N_270, N_272, 
        \state_ns_0_a2_1[0] , \state_ns_0_a2_0[0] , \state[7]_net_1 , 
        next_state_0_sqmuxa_1_1_a2_0_a2_0, \state_ns_i_0_0[2] , 
        un1_countlto15_13, un1_countlto15_5, un1_countlto15_4, 
        un1_countlto15_11, un1_countlto15_12, un1_countlto15_1, 
        un1_countlto15_0, un1_countlto15_9, un1_countlto15_7, 
        un1_countlto15_3, \state_RNO_1[5] , N_24, N_274, N_23, N_26, 
        next_state15_li, \state_RNIROJE[4]_net_1 , N_273, 
        \state[0]_net_1 , count_n7, count_n6, count_n5, count_n4, 
        count_n3, count_n2, count_n8, count_n9, count_n10, 
        \state_ns[7] , \state_ns[4] , \state[4]_net_1 , 
        \state_RNO_2[8] , count_n1, N_267, \state_ns[10] , 
        \state[12]_net_1 , \state_ns[12] , N_27, \state_ns[0] , 
        \state_ns[1] , \avg_count[1]_net_1 , \avg_count[0]_net_1 , 
        counte, \DWACT_ADD_CI_0_partial_sum[0] , I_10_2, 
        \DWACT_ADD_CI_0_TMP[0] , GND, VCC;
    
    DFN1E1C0 \count[5]  (.D(count_n5), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[5]_net_1 ));
    OA1A \state_RNO_0[0]  (.A(\state[10]_net_1 ), .B(N_33), .C(
        \state_ns_0_a2_8[0] ), .Y(\state_ns_0_a2_9[0] ));
    DFN1E1C0 \count[1]  (.D(count_n1), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[1]_net_1 ));
    OR2B \state_RNIBILG[4]  (.A(\state[4]_net_1 ), .B(
        \state[12]_net_1 ), .Y(N_273));
    DFN1E1C0 \count[10]  (.D(count_n10), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[10]_net_1 ));
    DFN1E1C0 \count[0]  (.D(N_267), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[0]_net_1 ));
    NOR2 \state_RNO_9[0]  (.A(calc_avg), .B(deriv_enable), .Y(
        \state_ns_0_a2_0[0] ));
    AOI1B \state_RNIOKMD4[10]  (.A(un1_countlto15_13), .B(
        un1_countlto15_12), .C(next_state_0_sqmuxa_1_1_a2_0_a2_0), .Y(
        N_62));
    DFN1C0 \state[13]  (.D(N_12), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_chg));
    DFN1E1C0 \count[14]  (.D(count_n14), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[14]_net_1 ));
    DFN1C0 \state[7]  (.D(\state_ns[7] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[7]_net_1 ));
    AX1C \count_RNO_0[14]  (.A(\count[13]_net_1 ), .B(count_c12), .C(
        \count[14]_net_1 ), .Y(count_n14_tz));
    OR2B \avg_count_RNIVG3T[1]  (.A(\avg_count[1]_net_1 ), .B(
        \avg_count[0]_net_1 ), .Y(next_state15_li));
    NOR2B \state_RNIROJE[4]  (.A(\state[4]_net_1 ), .B(avg_done), .Y(
        \state_RNIROJE[4]_net_1 ));
    DFN1C0 \state[5]  (.D(\state_RNO_1[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state_0[5] ));
    XA1B \count_RNO[7]  (.A(\count[7]_net_1 ), .B(count_c6), .C(N_62), 
        .Y(count_n7));
    AX1 \count_RNO[15]  (.A(N_62), .B(\count[15]_net_1 ), .C(N_94), .Y(
        count_n15));
    NOR3A \state_RNI6UI41[12]  (.A(\state[12]_net_1 ), .B(state_0_d0), 
        .C(state_0_0), .Y(N_12));
    NOR3C \count_RNI76NU1[7]  (.A(un1_countlto15_5), .B(
        un1_countlto15_4), .C(un1_countlto15_11), .Y(un1_countlto15_13)
        );
    NOR2B \count_RNITGCV2[12]  (.A(count_c11), .B(\count[12]_net_1 ), 
        .Y(count_c12));
    DFN1C0 \state[4]  (.D(\state_ns[4] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[4]_net_1 ));
    XA1B \count_RNO[2]  (.A(\count[2]_net_1 ), .B(count_c1), .C(N_62), 
        .Y(count_n2));
    NOR2B \count_RNI9U3L[2]  (.A(count_c1), .B(\count[2]_net_1 ), .Y(
        count_c2));
    NOR2 \count_RNI7L2E[1]  (.A(\count[2]_net_1 ), .B(\count[1]_net_1 )
        , .Y(un1_countlto15_1));
    AO1A \state_RNO[7]  (.A(N_46_1), .B(\state[7]_net_1 ), .C(calc_int)
        , .Y(\state_ns[7] ));
    DFN1C0 \state_1[2]  (.D(\state_RNI808O1[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable_1));
    NOR2A \state_RNO_0[5]  (.A(N_272), .B(\state[10]_net_1 ), .Y(N_24));
    DFN1C0 \state_0[2]  (.D(\state_RNI808O1[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable_0));
    XA1B \count_RNO[9]  (.A(count_c8), .B(\count[9]_net_1 ), .C(N_62), 
        .Y(count_n9));
    NOR2B \count_RNI8D2N2[11]  (.A(count_c10), .B(\count[11]_net_1 ), 
        .Y(count_c11));
    AO1 \state_RNIMF4H4[10]  (.A(sig_old_i_0), .B(sig_prev), .C(N_62), 
        .Y(counte));
    DFN1C0 \state[6]  (.D(int_enable), .CLK(clk_c), .CLR(n_rst_c), .Q(
        calc_int));
    NOR2 \state_RNO_6[0]  (.A(sum_enable), .B(\state[7]_net_1 ), .Y(
        \state_ns_0_a2_2[0] ));
    DFN1C0 \state[2]  (.D(\state_RNI808O1[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable));
    VCC VCC_i (.Y(VCC));
    XOR2 un1_avg_count_1_I_10 (.A(\avg_count[1]_net_1 ), .B(
        \DWACT_ADD_CI_0_TMP[0] ), .Y(I_10_2));
    NOR2 \count_RNIFT2E[5]  (.A(\count[6]_net_1 ), .B(\count[5]_net_1 )
        , .Y(un1_countlto15_3));
    XA1B \count_RNO[4]  (.A(\count[4]_net_1 ), .B(count_c3), .C(N_62), 
        .Y(count_n4));
    DFN1C0 \state[3]  (.D(avg_enable), .CLK(clk_c), .CLR(n_rst_c), .Q(
        calc_avg));
    NOR2B \count_RNI19E62[9]  (.A(count_c8), .B(\count[9]_net_1 ), .Y(
        count_c9));
    DFN1E1C0 \count[8]  (.D(count_n8), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[8]_net_1 ));
    XA1B \count_RNO[10]  (.A(count_c9), .B(\count[10]_net_1 ), .C(N_62)
        , .Y(count_n10));
    NOR2B \state_RNO[8]  (.A(\state[7]_net_1 ), .B(N_46_1), .Y(
        \state_RNO_2[8] ));
    NOR3B \state_RNO_1[0]  (.A(next_state15_li), .B(
        \state_RNIROJE[4]_net_1 ), .C(\state[10]_net_1 ), .Y(N_26));
    OR2A \state_RNIJHR3[7]  (.A(vd_rdy), .B(\state[7]_net_1 ), .Y(
        \state_ns_i_0_0[2] ));
    NOR2B \count_RNI5J2E[1]  (.A(\count[0]_net_1 ), .B(
        \count[1]_net_1 ), .Y(count_c1));
    DFN1E1C0 \count[15]  (.D(count_n15), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[15]_net_1 ));
    XA1B \count_RNO[3]  (.A(\count[3]_net_1 ), .B(count_c2), .C(N_62), 
        .Y(count_n3));
    NOR3 \state_RNI808O1[0]  (.A(N_274), .B(\state_ns_i_0_0[2] ), .C(
        N_23), .Y(\state_RNI808O1[0]_net_1 ));
    NOR2B \count_RNIKN631[4]  (.A(count_c3), .B(\count[4]_net_1 ), .Y(
        count_c4));
    DFN1E1C0 \count[11]  (.D(count_n11), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[11]_net_1 ));
    OA1 \state_RNO_0[12]  (.A(state_0_d0), .B(state_0_0), .C(
        \state[12]_net_1 ), .Y(N_27));
    DFN1C0 \state_0[13]  (.D(N_12), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_chg_0));
    XA1B \count_RNO[8]  (.A(count_c7), .B(\count[8]_net_1 ), .C(N_62), 
        .Y(count_n8));
    NOR3C \count_RNIRRJP1[1]  (.A(un1_countlto15_1), .B(
        un1_countlto15_0), .C(un1_countlto15_9), .Y(un1_countlto15_12));
    AO1A \state_RNO[10]  (.A(sum_rdy), .B(\state[10]_net_1 ), .C(
        sum_enable), .Y(\state_ns[10] ));
    DFN1E1C0 \count[13]  (.D(count_n13), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[13]_net_1 ));
    XA1B \count_RNO[5]  (.A(\count[5]_net_1 ), .B(count_c4), .C(N_62), 
        .Y(count_n5));
    XA1B \count_RNO[1]  (.A(\count[1]_net_1 ), .B(\count[0]_net_1 ), 
        .C(N_62), .Y(count_n1));
    XA1B \count_RNO[11]  (.A(count_c10), .B(\count[11]_net_1 ), .C(
        N_62), .Y(count_n11));
    NOR2 \count_RNIQFBF[15]  (.A(\count[15]_net_1 ), .B(
        \count[0]_net_1 ), .Y(un1_countlto15_0));
    NOR3B \state_RNO_4[0]  (.A(\state_ns_0_a2_2[0] ), .B(N_270), .C(
        N_272), .Y(\state_ns_0_a2_6[0] ));
    DFN1C0 \state[11]  (.D(N_62), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_enable));
    NOR2B \count_RNIR58A1[5]  (.A(count_c4), .B(\count[5]_net_1 ), .Y(
        count_c5));
    DFN1E1C0 \count[2]  (.D(count_n2), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[2]_net_1 ));
    DFN1P0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .PRE(n_rst_c), 
        .Q(\state[0]_net_1 ));
    NOR2B \count_RNIMMCV1[8]  (.A(count_c7), .B(\count[8]_net_1 ), .Y(
        count_c8));
    DFN1C0 \state[12]  (.D(\state_ns[12] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[12]_net_1 ));
    NOR2B \count_RNIEA5S[3]  (.A(count_c2), .B(\count[3]_net_1 ), .Y(
        count_c3));
    NOR2A \count_RNO_1[15]  (.A(\count[14]_net_1 ), .B(N_62), .Y(
        count_31_0));
    GND GND_i (.Y(GND));
    DFN1E1C0 \count[9]  (.D(count_n9), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[9]_net_1 ));
    NOR2B \state_RNIMIBL[10]  (.A(\state[10]_net_1 ), .B(sum_rdy), .Y(
        next_state_0_sqmuxa_1_1_a2_0_a2_0));
    XA1B \count_RNO[6]  (.A(\count[6]_net_1 ), .B(count_c5), .C(N_62), 
        .Y(count_n6));
    XA1B \count_RNO[12]  (.A(count_c11), .B(\count[12]_net_1 ), .C(
        N_62), .Y(count_n12));
    NOR2 \count_RNO[0]  (.A(\count[0]_net_1 ), .B(N_62), .Y(N_267));
    AND2 un1_avg_count_1_I_1 (.A(\avg_count[0]_net_1 ), .B(
        \state_RNIROJE[4]_net_1 ), .Y(\DWACT_ADD_CI_0_TMP[0] ));
    XOR2 un1_avg_count_1_I_8 (.A(\avg_count[0]_net_1 ), .B(
        \state_RNIROJE[4]_net_1 ), .Y(\DWACT_ADD_CI_0_partial_sum[0] ));
    NOR3B \state_RNO_5[0]  (.A(\state_ns_0_a2_1[0] ), .B(
        \state_ns_0_a2_0[0] ), .C(calc_error), .Y(\state_ns_0_a2_5[0] )
        );
    OR2 \state_RNIBILG_0[4]  (.A(\state[4]_net_1 ), .B(
        \state[12]_net_1 ), .Y(N_272));
    NOR2 \count_RNIJ13E[7]  (.A(\count[7]_net_1 ), .B(\count[8]_net_1 )
        , .Y(un1_countlto15_4));
    NOR3C \state_RNO_2[0]  (.A(un1_countlto15_12), .B(
        un1_countlto15_13), .C(sum_rdy), .Y(N_33));
    NOR2 \count_RNIUJBF[9]  (.A(\count[9]_net_1 ), .B(
        \count[10]_net_1 ), .Y(un1_countlto15_5));
    NOR2B \count_RNIKAOE2[10]  (.A(count_c9), .B(\count[10]_net_1 ), 
        .Y(count_c10));
    AO1A \state_RNO[4]  (.A(avg_done), .B(\state[4]_net_1 ), .C(
        calc_avg), .Y(\state_ns[4] ));
    DFN1E1C0 \count[6]  (.D(count_n6), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[6]_net_1 ));
    OR2 \state_RNO[12]  (.A(N_27), .B(pwm_enable), .Y(\state_ns[12] ));
    DFN1C0 \state[10]  (.D(\state_ns[10] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[10]_net_1 ));
    DFN1E1C0 \count[3]  (.D(count_n3), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[3]_net_1 ));
    DFN1C0 \state[1]  (.D(\state_ns[1] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(calc_error));
    NOR2 \state_RNO_8[0]  (.A(pwm_enable), .B(calc_int), .Y(
        \state_ns_0_a2_1[0] ));
    DFN1C0 \state[8]  (.D(\state_RNO_2[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(deriv_enable));
    NOR2B \count_RNIC5BO1[7]  (.A(count_c6), .B(\count[7]_net_1 ), .Y(
        count_c7));
    NOR3A \state_RNO[5]  (.A(calc_error), .B(\state[7]_net_1 ), .C(
        N_24), .Y(\state_RNO_1[5] ));
    NOR2 \count_RNIDAKG[14]  (.A(\count[14]_net_1 ), .B(
        \count[13]_net_1 ), .Y(un1_countlto15_7));
    CLKINT \state_RNIV2C2[5]  (.A(\state_0[5] ), .Y(int_enable));
    NOR2A \count_RNO[14]  (.A(count_n14_tz), .B(N_62), .Y(count_n14));
    NOR3A \count_RNIMG811[11]  (.A(un1_countlto15_7), .B(
        \count[12]_net_1 ), .C(\count[11]_net_1 ), .Y(
        un1_countlto15_11));
    NOR3A \count_RNIQM5S[3]  (.A(un1_countlto15_3), .B(
        \count[3]_net_1 ), .C(\count[4]_net_1 ), .Y(un1_countlto15_9));
    XA1B \count_RNO[13]  (.A(count_c12), .B(\count[13]_net_1 ), .C(
        N_62), .Y(count_n13));
    DFN1C0 \state[9]  (.D(deriv_enable), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(sum_enable));
    NOR3A \state_RNIGUA11[0]  (.A(N_273), .B(\state[10]_net_1 ), .C(
        \state[0]_net_1 ), .Y(N_274));
    DFN1C0 \avg_count[0]  (.D(\DWACT_ADD_CI_0_partial_sum[0] ), .CLK(
        clk_c), .CLR(n_rst_c), .Q(\avg_count[0]_net_1 ));
    OR2B \state_RNO_7[0]  (.A(vd_rdy), .B(\state[0]_net_1 ), .Y(N_270));
    NOR2B \count_RNI3L9H1[6]  (.A(count_c5), .B(\count[6]_net_1 ), .Y(
        count_c6));
    AO1A \state_RNO[0]  (.A(int_enable), .B(\state_ns_0_a2_9[0] ), .C(
        N_26), .Y(\state_ns[0] ));
    DFN1C0 \avg_count[1]  (.D(I_10_2), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \avg_count[1]_net_1 ));
    NOR3C \count_RNO_0[15]  (.A(\count[13]_net_1 ), .B(count_c12), .C(
        count_31_0), .Y(N_94));
    NOR3B \state_RNO_3[0]  (.A(\state_ns_0_a2_6[0] ), .B(
        \state_ns_0_a2_5[0] ), .C(avg_enable), .Y(\state_ns_0_a2_8[0] )
        );
    DFN1E1C0 \count[4]  (.D(count_n4), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[4]_net_1 ));
    DFN1E1C0 \count[12]  (.D(count_n12), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[12]_net_1 ));
    NOR2A \state_RNO[1]  (.A(\state_RNIROJE[4]_net_1 ), .B(
        next_state15_li), .Y(\state_ns[1] ));
    NOR2 \state_RNI5G1J[0]  (.A(\state[0]_net_1 ), .B(N_272), .Y(N_23));
    DFN1E1C0 \count[7]  (.D(count_n7), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[7]_net_1 ));
    
endmodule


module sig_gen_6(
       primary_5_c,
       n_rst_c,
       clk_c,
       sig_old_i_0,
       sig_prev
    );
input  primary_5_c;
input  n_rst_c;
input  clk_c;
output sig_old_i_0;
output sig_prev;

    wire sig_prev_i, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(clk_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev_inst_1 (.D(primary_5_c), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(sig_prev));
    INV sig_old_RNO (.A(sig_prev), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module pid_sum_13s_4_2(
       integral_i,
       integral,
       sr_new,
       integral_1_0,
       sr_new_1_0,
       sr_new_0_0,
       derivative_0,
       integral_0_0,
       sum_39,
       sum_14,
       sum_19,
       sum_20,
       sum_22,
       sum_13,
       sum_17,
       sum_18,
       sum_23,
       sum_21,
       sum_16,
       sum_15,
       sum_12,
       sum_11,
       sum_6,
       sum_10,
       sum_9,
       sum_5,
       sum_8,
       sum_7,
       sum_4,
       sum_2_d0,
       sum_1_d0,
       sum_0_d0,
       sum_3,
       sum_0_0,
       sum_1_0,
       sum_2_0,
       sum_enable,
       sum_rdy,
       n_rst_c,
       clk_c
    );
input  [25:24] integral_i;
input  [25:6] integral;
input  [12:0] sr_new;
input  integral_1_0;
input  sr_new_1_0;
input  sr_new_0_0;
input  derivative_0;
input  integral_0_0;
output sum_39;
output sum_14;
output sum_19;
output sum_20;
output sum_22;
output sum_13;
output sum_17;
output sum_18;
output sum_23;
output sum_21;
output sum_16;
output sum_15;
output sum_12;
output sum_11;
output sum_6;
output sum_10;
output sum_9;
output sum_5;
output sum_8;
output sum_7;
output sum_4;
output sum_2_d0;
output sum_1_d0;
output sum_0_d0;
output sum_3;
output sum_0_0;
output sum_1_0;
output sum_2_0;
input  sum_enable;
output sum_rdy;
input  n_rst_c;
input  clk_c;

    wire \next_sum[39] , N_416, \state_0[1]_net_1 , 
        \state_RNIEBE9[0]_net_1 , \state_2[2]_net_1 , 
        \state_1[2]_net_1 , \state_0[2]_net_1 , \state_0[3]_net_1 , 
        \state[6]_net_1 , N_416_0, \un1_next_sum_1_iv_0[26] , 
        \un1_next_sum_0_iv_0[25] , next_sum_1_sqmuxa, N_12, N_10, 
        \DWACT_FINC_E[0] , N_5, \DWACT_FINC_E[4] , N_2, 
        \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , N_25, N_23, 
        \DWACT_FINC_E_0[0] , N_18, \DWACT_FINC_E_0[4] , N_15, 
        \DWACT_FINC_E_0[7] , \DWACT_FINC_E_0[6] , 
        ADD_40x40_fast_I448_Y_0, \sumreg[30]_net_1 , 
        \un1_next_sum_1_iv[26] , ADD_40x40_fast_I447_Y_0, 
        \sumreg[29]_net_1 , ADD_40x40_fast_I456_Y_0, 
        \sumreg[38]_net_1 , ADD_40x40_fast_I449_Y_0, 
        \sumreg[31]_net_1 , ADD_40x40_fast_I453_Y_0, 
        \sumreg[35]_net_1 , ADD_40x40_fast_I454_Y_0, 
        \sumreg[36]_net_1 , ADD_40x40_fast_I455_Y_0, 
        \sumreg[37]_net_1 , ADD_40x40_fast_I451_Y_0, 
        \sumreg[33]_net_1 , ADD_40x40_fast_I452_Y_0, 
        \sumreg[34]_net_1 , ADD_40x40_fast_I347_Y_0, N787, N772, N771, 
        ADD_40x40_fast_I457_Y_0, ADD_40x40_fast_I446_Y_0, 
        \sumreg[28]_net_1 , ADD_40x40_fast_I450_Y_0, 
        \sumreg[32]_net_1 , ADD_40x40_fast_I379_Y_4, I268_un1_Y, 
        ADD_40x40_fast_I379_Y_2, I332_un1_Y, N596, 
        ADD_40x40_fast_I379_Y_0, N681, ADD_40x40_fast_I346_Y_0, N785, 
        N770, N769, ADD_40x40_fast_I382_Y_1, N762, N777, 
        ADD_40x40_fast_I382_Y_0, N679, N687, ADD_40x40_fast_I381_Y_2, 
        N760, N775, ADD_40x40_fast_I381_Y_1, N600, N685, 
        ADD_40x40_fast_I445_Y_0, \sumreg[27]_net_1 , 
        ADD_40x40_fast_I432_Y_0, \un1_next_sum[14] , 
        ADD_40x40_fast_I380_Y_2, N758, N773, ADD_40x40_fast_I380_Y_1, 
        N598, N594, N683, ADD_40x40_fast_I437_Y_0, \un1_next_sum[19] , 
        ADD_40x40_fast_I438_Y_0, \un1_next_sum_2[4] , 
        \un1_next_sum_iv_0[20] , ADD_40x40_fast_I383_Y_1, N764, N779, 
        ADD_40x40_fast_I383_Y_0, N689, ADD_40x40_fast_I384_Y_2, 
        ADD_40x40_fast_I384_Y_0, I278_un1_Y, I384_un1_Y, N691, N684, 
        ADD_40x40_fast_I444_Y_0, \sumreg[26]_net_1 , 
        ADD_40x40_fast_I443_Y_0, \sumreg[25]_net_1 , 
        \un1_next_sum_0_iv[25] , ADD_40x40_fast_I440_Y_0, 
        \un1_next_sum_iv_0[22] , ADD_40x40_fast_I378_Y_3, N754, 
        ADD_40x40_fast_I378_Y_2, ADD_40x40_fast_I378_Y_0, 
        ADD_40x40_fast_I385_Y_1, N768, N783, ADD_40x40_fast_I385_Y_0, 
        N693, N686, ADD_40x40_fast_I431_Y_0, \un1_next_sum[13] , 
        ADD_40x40_fast_I442_Y_0, \un1_next_sum_iv_0[24] , 
        \sumreg[24]_net_1 , ADD_40x40_fast_I435_Y_0, 
        \un1_next_sum[17] , ADD_40x40_fast_I436_Y_0, 
        \un1_next_sum_iv_1[18] , \un1_next_sum_iv_2[18] , 
        ADD_40x40_fast_I441_Y_0, \un1_next_sum_iv_0[23] , 
        ADD_40x40_fast_I439_Y_0, \un1_next_sum[21] , 
        ADD_40x40_fast_I434_Y_0, \un1_next_sum_iv_1[16] , 
        \un1_next_sum_iv_2[16] , ADD_40x40_fast_I433_Y_0, 
        \un1_next_sum[15] , ADD_40x40_fast_I346_un1_Y_0, N786, 
        ADD_40x40_fast_I430_Y_0, \un1_next_sum[12] , 
        ADD_40x40_fast_I352_Y_0, N797, N782, N781, 
        ADD_40x40_fast_I353_Y_0, N799, N784, 
        ADD_40x40_fast_I379_un1_Y_0, N756, N872, 
        ADD_40x40_fast_I429_Y_0, \un1_next_sum[11] , 
        ADD_40x40_fast_I380_un1_Y_0, N874, N821, 
        ADD_40x40_fast_I424_Y_0, \un1_next_sum[6] , 
        ADD_40x40_fast_I428_Y_0, \un1_next_sum[10] , 
        ADD_40x40_fast_I427_Y_0, \un1_next_sum_iv_1[9] , 
        \un1_next_sum_iv_2[9] , ADD_40x40_fast_I378_un1_Y_0, N870, 
        N817, ADD_40x40_fast_I352_un1_Y_0, N798, 
        ADD_40x40_fast_I423_Y_0, \un1_next_sum_iv_0[5] , 
        ADD_40x40_fast_I426_Y_0, \un1_next_sum[8] , 
        ADD_40x40_fast_I353_un1_Y_0, N800, ADD_40x40_fast_I425_Y_0, 
        \un1_next_sum_iv_1[7] , \un1_next_sum_iv_2[7] , 
        ADD_40x40_fast_I422_Y_0, \un1_next_sum_iv_0[4] , 
        ADD_40x40_fast_I420_Y_0, \un1_next_sum[0] , 
        ADD_40x40_fast_I419_Y_0, ADD_40x40_fast_I257_Y_1, N475, N472, 
        N661, ADD_40x40_fast_I201_Y_0, N601, N597, 
        ADD_40x40_fast_I195_Y_0, ADD_40x40_fast_I197_Y_0, 
        ADD_40x40_fast_I187_Y_0, ADD_22x22_fast_I176_Y_0, 
        \i_adj[16]_net_1 , \i_adj[18]_net_1 , ADD_22x22_fast_I126_Y_1, 
        N371, N378, ADD_22x22_fast_I126_Y_0, N335, N332, N331, 
        ADD_22x22_fast_I142_Y_0_1, ADD_22x22_fast_I142_Y_0_a3_0, N329, 
        ADD_22x22_fast_I142_Y_0_0, \i_adj[20]_net_1 , N_7, 
        ADD_22x22_fast_I168_Y_0, \i_adj[10]_net_1 , \i_adj[8]_net_1 , 
        ADD_22x22_fast_I126_un1_Y_0, N379, 
        ADD_22x22_fast_I142_Y_0_a3_1, N330, ADD_40x40_fast_I418_Y_0, 
        ADD_22x22_fast_I177_Y_0, \i_adj[19]_net_1 , \i_adj[17]_net_1 , 
        ADD_22x22_fast_I130_Y_0, N386, ADD_40x40_fast_I421_Y_0, N743, 
        ADD_22x22_fast_I142_Y_0_o3_0_0, N337, N334, N333, 
        ADD_22x22_fast_I128_Y_0, N382, N375, N374, 
        ADD_22x22_fast_I164_Y_0, \i_adj[4]_net_1 , \i_adj[6]_net_1 , 
        ADD_22x22_fast_I143_Y_2, N367, ADD_22x22_fast_I143_Y_1, N328, 
        ADD_22x22_fast_I143_Y_0, N314, ADD_22x22_fast_I144_Y_2, 
        ADD_22x22_fast_I144_un1_Y_0, N425, ADD_22x22_fast_I144_Y_1, 
        N369, N376, ADD_22x22_fast_I144_Y_0, 
        ADD_22x22_fast_I130_un1_Y_0, N387, \un1_next_sum_iv_0[21] , 
        \ireg[21]_net_1 , \ireg[20]_net_1 , \un1_next_sum_iv_0[19] , 
        \ireg[19]_net_1 , \ireg[23]_net_1 , \ireg[24]_net_1 , 
        \ireg[5]_net_1 , \ireg[22]_net_1 , \ireg[4]_net_1 , 
        ADD_22x22_fast_I170_Y_0, \i_adj[12]_net_1 , 
        ADD_22x22_fast_I169_Y_0, \i_adj[9]_net_1 , \i_adj[11]_net_1 , 
        \un24_next_sum_m[16] , next_sum_0_sqmuxa_1, 
        \un3_next_sum_m[16] , \ireg[16]_net_1 , \preg_m[16] , 
        \un1_next_sum_iv_2[13] , \un24_next_sum_m[13] , 
        \un3_next_sum_m[13] , \un1_next_sum_iv_1[13] , 
        \preg[13]_net_1 , next_sum_1_sqmuxa_2, \ireg_m[13] , 
        \un1_next_sum_iv_2[11] , \un24_next_sum_m[11] , 
        \un3_next_sum_m[11] , \un1_next_sum_iv_1[11] , 
        \preg[11]_net_1 , \ireg_m[11] , \un1_next_sum_iv_2[17] , 
        \un3_next_sum_m[17] , \un1_next_sum_iv_0[17] , 
        \un1_next_sum_iv_1[17] , \ireg[17]_net_1 , \preg_m[17] , 
        \un24_next_sum_m[17] , \un1_next_sum_iv_2[8] , 
        \un3_next_sum_m[8] , \un1_next_sum_iv_0[8] , 
        \un1_next_sum_iv_1[8] , \preg[8]_net_1 , \ireg_m[8] , 
        \un24_next_sum_m[8] , \un24_next_sum_m[18] , 
        \un3_next_sum_m[18] , \ireg[18]_net_1 , \preg_m[18] , 
        \un1_next_sum_iv_2[15] , \un24_next_sum_m[15] , 
        \un3_next_sum_m[15] , \un1_next_sum_iv_1[15] , 
        \ireg[15]_net_1 , \preg_m[15] , \un24_next_sum_m[7] , 
        \un3_next_sum_m[7] , \preg[7]_net_1 , \ireg_m[7] , 
        \un1_next_sum_iv_2[10] , \un3_next_sum_m[10] , 
        \un1_next_sum_iv_0[10] , \un1_next_sum_iv_1[10] , 
        \preg[10]_net_1 , \ireg_m[10] , \un24_next_sum_m[10] , 
        \un1_next_sum_iv_2[6] , \un3_next_sum_m[6] , 
        \un1_next_sum_iv_0[6] , \un1_next_sum_iv_1[6] , 
        \preg[6]_net_1 , \ireg_m[6] , \un24_next_sum_m[6] , 
        \un1_next_sum_iv_2[14] , \un24_next_sum_m[14] , 
        \un3_next_sum_m[14] , \un1_next_sum_iv_1[14] , 
        \ireg[14]_net_1 , \preg_m[14] , \un1_next_sum_iv_2[12] , 
        \ireg[12]_net_1 , next_sum_0_sqmuxa, \un1_next_sum_iv_0[12] , 
        \un1_next_sum_iv_1[12] , \preg[12]_net_1 , \ireg_m[12] , 
        \un24_next_sum_m[12] , \un24_next_sum_m[9] , 
        \un3_next_sum_m[9] , \preg[9]_net_1 , \ireg_m[9] , 
        next_sum_0_sqmuxa_2, ADD_22x22_fast_I128_un1_Y_0, N383, 
        ADD_22x22_fast_I142_Y_0_a3_3_0, N338, \state[4]_net_1 , 
        ADD_22x22_fast_I129_Y_0, N384, N377, ADD_22x22_fast_I131_Y_0, 
        N345, N342, N341, ADD_22x22_fast_I165_Y_0, \i_adj[5]_net_1 , 
        \i_adj[7]_net_1 , ADD_22x22_fast_I129_un1_Y_0, N385, N266, 
        ADD_22x22_fast_I162_Y_0, \i_adj[2]_net_1 , 
        ADD_22x22_fast_I163_Y_0, \i_adj[3]_net_1 , N_9, 
        ADD_m8_i_a4_0_0, ADD_m8_i_o4_1, ADD_m8_i_a4_0, ADD_m8_i_a4, 
        N_232, N492, N_11, I143_un1_Y, N407, N423, N359, N494, 
        I122_un1_Y, I126_un1_Y, I112_un1_Y, N504, N528, 
        \next_ireg_3[12] , \next_ireg_3[24] , \next_ireg_3[22] , 
        \next_ireg_3[20] , \i_adj[14]_net_1 , \next_ireg_3[25] , 
        \i_adj[21]_net_1 , \next_ireg_3[17] , \i_adj[13]_net_1 , N513, 
        N816, N734, N682, I378_un1_Y, N1021, I330_un1_Y, N1049, 
        I290_un1_Y, I350_un1_Y, N778, N794, N1097, N1029, I382_un1_Y, 
        I338_un1_Y, N878, N846, N595, N680, N1058, N1106, 
        \un3_next_sum_m[25] , \ireg_m[25] , \next_ireg_3[13] , N525, 
        \next_ireg_3[11] , N531, \next_ireg_3[9] , N396, I131_un1_Y, 
        I106_un1_Y, N389, N381, \state[1]_net_1 , \state[5]_net_1 , 
        \next_ireg_3[7] , \i_adj[1]_net_1 , I348_un1_Y, N774, N790, 
        N1091, N1043, I286_un1_Y, N1055, N1103, I380_un1_Y, N1025, 
        I334_un1_Y, I381_un1_Y, N876, N823, N844, N1027, I336_un1_Y, 
        N882, N666, N850, N1033, N881, I385_un1_Y, N884, N852, N1035, 
        I344_un1_Y, N1037, N1085, \next_ireg_3[8] , \next_ireg_3[10] , 
        N394, \next_ireg_3[16] , N422, I132_un1_Y, \next_ireg_3[15] , 
        N424, I133_un1_Y, \next_ireg_3[19] , \i_adj[15]_net_1 , N507, 
        \next_ireg_3[21] , \next_ireg_3[23] , I124_un1_Y, 
        \next_ireg_3[18] , N510, \next_ireg_3[14] , N1031, I383_un1_Y, 
        I340_un1_Y, N880, N745, N848, N1023, N819, N1052, I292_un1_Y, 
        I351_un1_Y, N780, N796, N1100, N1046, I288_un1_Y, I349_un1_Y, 
        N776, N792, N1094, N1040, I347_un1_Y, N788, N1088, N599, N740, 
        N484, N481, \next_sum[4] , \state[2]_net_1 , \next_sum[5] , 
        \next_sum[7] , \next_sum[10] , \next_sum[11] , \next_sum[12] , 
        \next_sum[13] , \next_sum[14] , \next_sum[17] , N1079, 
        \next_sum[18] , N1076, \next_sum[19] , N1073, \next_sum[20] , 
        N1070, \next_sum[21] , N1067, \next_sum[22] , N1064, 
        \next_sum[26] , \next_sum[30] , \next_sum[34] , \next_sum[38] , 
        N272, N278, N279, N284, N288, N290, N291, N294, N343, N293, 
        N347, N287, N355, N344, N354, N350, N282, N348, N346, N340, 
        N300, N339, N296, N299, N275, \i_adj[0]_net_1 , N388, N353, 
        N349, \next_ireg_3[6] , N357, N269, N273, N281, N722, N645, 
        N641, N791, N717, N710, N709, N718, N714, N804, N730, N811, 
        N737, N729, N812, N738, N879, N795, N721, N713, N636, N633, 
        N632, N519, N520, N637, N514, N698, N706, N625, N629, N526, 
        N640, N513_0, N628, N525_0, N644, N501, N505, N504_0, N507_0, 
        N510_0, N511, N638, N639, N642, N643, N716, N635, N732, N651, 
        N655, I186_un1_Y, N662, N739, N658, N806, N724, N813, N731, 
        N814, I260_un1_Y, N712, N631, N711, N634, N630, N522, N528_0, 
        N531_0, N532, N534, N540, N541, N606, N623, N538, N624, N626, 
        N627, N516, N700, N619, N705, N707, N708, N715, N692, N697, 
        I222_un1_Y, N699, N789, N723, N803, N805, N871, N873, N875, 
        N807, N808, N877, \inf_abs1_5[0] , \inf_abs1_5[1] , 
        \inf_abs1_a_2[1] , \inf_abs1_5[2] , \inf_abs1_a_2[2] , 
        \inf_abs1_5[3] , \inf_abs1_a_2[3] , \inf_abs1_5[4] , 
        \inf_abs1_a_2[4] , \inf_abs1_5[5] , \inf_abs1_a_2[5] , 
        \inf_abs1_5[7] , \inf_abs1_a_2[7] , \inf_abs1_5[8] , 
        \inf_abs1_a_2[8] , \inf_abs1_5[9] , \inf_abs1_a_2[9] , 
        \inf_abs1_5[10] , \inf_abs1_a_2[10] , \inf_abs2_5[0] , 
        \inf_abs2_5[1] , \inf_abs2_a_0[1] , \inf_abs2_5[2] , 
        \inf_abs2_a_0[2] , \inf_abs2_5[4] , \inf_abs2_a_0[4] , 
        \inf_abs2_5[5] , \inf_abs2_a_0[5] , \inf_abs2_5[6] , 
        \inf_abs2_a_0[6] , \inf_abs2_5[8] , \inf_abs2_a_0[8] , 
        \inf_abs2_5[9] , \inf_abs2_a_0[9] , \inf_abs2_5[10] , 
        \inf_abs2_a_0[10] , \inf_abs2_5[11] , \inf_abs2_a_0[11] , 
        \inf_abs2_5[12] , \inf_abs2_a_0[12] , \inf_abs2_5[13] , 
        \inf_abs2_a_0[13] , \inf_abs2_5[14] , \inf_abs2_a_0[14] , 
        \inf_abs2_5[15] , \inf_abs2_a_0[15] , \inf_abs2_5[16] , 
        \inf_abs2_a_0[16] , \inf_abs1_5[12] , \inf_abs1_a_2[12] , 
        \state[3]_net_1 , \ireg[6]_net_1 , \ireg[7]_net_1 , 
        \ireg[10]_net_1 , \ireg[11]_net_1 , \preg[14]_net_1 , 
        \preg[17]_net_1 , \preg[18]_net_1 , N704, N703, N622, N537, 
        \next_sum[31] , \next_sum[28] , \next_sum[27] , \next_sum[23] , 
        N1061, N883, N1082, I361_un1_Y, \next_sum[32] , \next_sum[16] , 
        N609, \next_sum[36] , \next_sum[33] , I214_un1_Y, N610, N608, 
        N607, \next_sum[37] , \next_sum[25] , \preg[15]_net_1 , 
        \inf_abs1_5[11] , \inf_abs1_a_2[11] , N_228, \preg[16]_net_1 , 
        \ireg[13]_net_1 , N358, N270, I87_un1_Y, N356, \state_ns[0] , 
        N688, N611, I138_un1_Y, N614, N615, N694, N701, N702, N613, 
        N617, N550, N616, N612, N620, N549, I218_un1_Y, N695, 
        \ireg[25]_net_1 , N618, I142_un1_Y, N544, N543, I64_un1_Y, 
        N621, I115_un1_Y, N392, N393, \next_sum[24] , \next_sum[29] , 
        \next_sum[35] , N602, N603, N793, N604, N605, N690, N802, N869, 
        N801, I318_un1_Y, N809, N728, N736, N735, N727, N720, N719, 
        N654, N650, N647, N646, N471, N664, I116_un1_Y, N741, N660, 
        \next_sum[9] , \next_sum[1] , \next_sum[2] , \next_sum[3] , 
        N726, N815, N733, I321_un1_Y, N480, N483, I108_un1_Y, 
        \ireg[9]_net_1 , \ireg[8]_net_1 , N495, N498, N487, N486, N493, 
        N492_0, N499, N489, N648, N649, N652, N657, N656, N653, N725, 
        \next_sum[8] , \next_sum[6] , \next_sum[0] , \inf_abs2_5[3] , 
        \inf_abs2_a_0[3] , \inf_abs1_5[6] , \inf_abs1_a_2[6] , 
        \inf_abs2_5[7] , \inf_abs2_a_0[7] , \inf_abs2_5[21] , 
        \inf_abs2_a_0[21] , \inf_abs2_5[20] , \inf_abs2_a_0[20] , 
        \inf_abs2_5[19] , \inf_abs2_a_0[19] , \inf_abs2_5[18] , 
        \inf_abs2_a_0[18] , \inf_abs2_5[17] , \inf_abs2_a_0[17] , N336, 
        N306, N302, N305, N312, N308, N311, N391, N390, I86_un1_Y, 
        N352, N351, \next_sum[15] , \p_adj[0]_net_1 , \p_adj[1]_net_1 , 
        \p_adj[2]_net_1 , \p_adj[3]_net_1 , \p_adj[4]_net_1 , 
        \p_adj[5]_net_1 , \p_adj[6]_net_1 , \p_adj[7]_net_1 , 
        \p_adj[8]_net_1 , \p_adj[9]_net_1 , \p_adj[10]_net_1 , 
        \p_adj[11]_net_1 , \p_adj[12]_net_1 , N_6, \DWACT_FINC_E[28] , 
        \DWACT_FINC_E[13] , \DWACT_FINC_E[15] , N_7_0, 
        \DWACT_FINC_E[14] , N_8, \DWACT_FINC_E[9] , \DWACT_FINC_E[12] , 
        N_9_0, \DWACT_FINC_E[10] , \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[5] , N_10_0, \DWACT_FINC_E[11] , N_11_0, N_12_0, 
        N_13, \DWACT_FINC_E[8] , N_14, N_16, N_17, \DWACT_FINC_E[3] , 
        N_19, N_20, N_21, \DWACT_FINC_E[1] , N_22, N_24, N_3, 
        \DWACT_FINC_E_0[2] , \DWACT_FINC_E_0[5] , N_4, 
        \DWACT_FINC_E_0[3] , N_6_0, N_7_1, N_8_0, \DWACT_FINC_E_0[1] , 
        N_9_1, N_11_1, GND, VCC;
    
    DFN1E1C0 \sumreg[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(sum_39));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I77_Y (.A(sum_19), .B(
        \un1_next_sum[19] ), .C(N532), .Y(N627));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_o3_0 (.A(
        ADD_22x22_fast_I142_Y_0_a3_3_0), .B(N513), .C(
        ADD_22x22_fast_I142_Y_0_o3_0_0), .Y(N_11));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I19_G0N (.A(\un1_next_sum[19] )
        , .B(sum_19), .Y(N528_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I14_P0N (.A(\un1_next_sum[14] ), 
        .B(sum_14), .Y(N514));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I46_Y (.A(\sumreg[34]_net_1 ), 
        .B(\sumreg[35]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N596)
        );
    XA1B \sumreg_RNO[10]  (.A(N1100), .B(ADD_40x40_fast_I428_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[10] ));
    MX2 \p_adj_RNO[2]  (.A(sr_new[2]), .B(\inf_abs1_a_2[2] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[2] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I336_un1_Y (.A(N844), .B(N875), 
        .Y(I336_un1_Y));
    XA1B \sumreg_RNO[11]  (.A(N1097), .B(ADD_40x40_fast_I429_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[11] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_0 (.A(N333), .B(N330), .C(
        N329), .Y(ADD_22x22_fast_I144_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I241_Y (.A(N726), .B(N718), .Y(
        N800));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I114_Y (.A(N471), .B(
        \un1_next_sum[0] ), .C(sum_1_d0), .Y(N664));
    DFN1E1C0 \i_adj[19]  (.D(\inf_abs2_5[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[19]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I113_Y (.A(N389), .B(N396), .C(
        N388), .Y(N525));
    DFN1E1C0 \sumreg[23]  (.D(\next_sum[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_23));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I290_un1_Y (.A(N793), .B(N778), 
        .Y(I290_un1_Y));
    XA1 \ireg_RNIHAEP[21]  (.A(integral_0_0), .B(\ireg[21]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[21] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I128_un1_Y_0 (.A(N383), .B(N375)
        , .Y(ADD_22x22_fast_I128_un1_Y_0));
    NOR3B inf_abs1_a_2_I_19 (.A(\DWACT_FINC_E_0[2] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[6]), .Y(N_7_1));
    OA1 next_ireg_3_0_ADD_22x22_fast_I33_Y (.A(\i_adj[12]_net_1 ), .B(
        \i_adj[14]_net_1 ), .C(N300), .Y(N338));
    AND3 inf_abs2_a_0_I_30 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E_0[6] ));
    MX2 \i_adj_RNO[5]  (.A(integral[11]), .B(\inf_abs2_a_0[5] ), .S(
        integral_1_0), .Y(\inf_abs2_5[5] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I304_Y (.A(N807), .B(N792), .C(
        N791), .Y(N875));
    DFN1E1C0 \sumreg[38]  (.D(\next_sum[38] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[38]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I126_un1_Y_0 (.A(N371), .B(N379)
        , .Y(ADD_22x22_fast_I126_un1_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I361_Y (.A(I361_un1_Y), .B(N883), 
        .Y(N1082));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I201_Y_0 (.A(N601), .B(N597), 
        .Y(ADD_40x40_fast_I201_Y_0));
    DFN1E1C0 \sumreg[5]  (.D(\next_sum[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416), .Q(sum_5));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I248_Y (.A(N733), .B(N726), .C(
        N725), .Y(N807));
    DFN1E1C0 \sumreg[20]  (.D(\next_sum[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_20));
    NOR3B \preg_RNI8RBI[14]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[14]_net_1 ), .Y(\un24_next_sum_m[14] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I128_Y (.A(
        ADD_22x22_fast_I128_un1_Y_0), .B(N528), .C(
        ADD_22x22_fast_I128_Y_0), .Y(N504));
    NOR2 inf_abs2_a_0_I_57 (.A(integral[24]), .B(integral[25]), .Y(
        \DWACT_FINC_E[14] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I347_Y_0 (.A(N787), .B(N772), .C(
        N771), .Y(ADD_40x40_fast_I347_Y_0));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I52_Y (.A(\sumreg[31]_net_1 ), 
        .B(\sumreg[32]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N602)
        );
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I199_Y (.A(N599), .B(N595), .C(
        N684), .Y(N758));
    DFN1E1C0 \sumreg[13]  (.D(\next_sum[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_13));
    NOR3B \ireg_RNIIADP[13]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[13]_net_1 ), .Y(\un3_next_sum_m[13] ));
    OR2 \preg_RNIA9581[8]  (.A(next_sum_0_sqmuxa_1), .B(
        \un24_next_sum_m[8] ), .Y(\un1_next_sum_iv_0[8] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I354_Y (.A(N870), .B(N817), .C(
        N869), .Y(N1061));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I214_Y (.A(I214_un1_Y), .B(N691), 
        .Y(N773));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I353_un1_Y_0 (.A(N800), .B(
        N784), .Y(ADD_40x40_fast_I353_un1_Y_0));
    DFN1E1C0 \i_adj[2]  (.D(\inf_abs2_5[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[2]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I225_Y (.A(N702), .B(N710), .Y(
        N784));
    NOR3A inf_abs1_a_2_I_13 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .C(
        sr_new[4]), .Y(N_9_1));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I436_Y_0 (.A(
        \un1_next_sum_iv_1[18] ), .B(\un1_next_sum_iv_2[18] ), .C(
        sum_18), .Y(ADD_40x40_fast_I436_Y_0));
    DFN1E1C0 \sumreg[27]  (.D(\next_sum[27] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[27]_net_1 ));
    DFN1E1C0 \sumreg[10]  (.D(\next_sum[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_10));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I381_Y_2 (.A(N760), .B(N775), .C(
        ADD_40x40_fast_I381_Y_1), .Y(ADD_40x40_fast_I381_Y_2));
    OR2 next_ireg_3_0_ADD_22x22_fast_I15_P0N (.A(\i_adj[17]_net_1 ), 
        .B(\i_adj[15]_net_1 ), .Y(N312));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I308_Y (.A(N811), .B(N796), .C(
        N795), .Y(N879));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I444_Y_0 (.A(
        \sumreg[26]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I444_Y_0));
    XA1B \sumreg_RNO[22]  (.A(N1064), .B(ADD_40x40_fast_I440_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[22] ));
    OR2 \state_RNI9CV41[4]  (.A(\un1_next_sum_0_iv_0[25] ), .B(
        next_sum_1_sqmuxa), .Y(\un1_next_sum_1_iv_0[26] ));
    OR2 \ireg_RNIKURG3[17]  (.A(\un1_next_sum_iv_2[17] ), .B(
        \un1_next_sum_iv_1[17] ), .Y(\un1_next_sum[17] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I171_Y (.A(N647), .B(N643), .Y(
        N724));
    OR2 next_ireg_3_0_ADD_22x22_fast_I11_P0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(N300));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I443_Y_0 (.A(
        \sumreg[25]_net_1 ), .B(\un1_next_sum_0_iv[25] ), .Y(
        ADD_40x40_fast_I443_Y_0));
    AND2 inf_abs2_a_0_I_44 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E[9] ), .Y(\DWACT_FINC_E[10] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I18_P0N (.A(
        \un1_next_sum_iv_1[18] ), .B(\un1_next_sum_iv_2[18] ), .C(
        sum_18), .Y(N526));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I166_Y (.A(N642), .B(N639), .C(
        N638), .Y(N719));
    OA1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_0_0 (.A(
        \i_adj[18]_net_1 ), .B(\i_adj[20]_net_1 ), .C(N_9), .Y(
        ADD_22x22_fast_I142_Y_0_a3_0));
    AX1D next_ireg_3_0_ADD_22x22_fast_I168_Y (.A(N386), .B(I112_un1_Y), 
        .C(ADD_22x22_fast_I168_Y_0), .Y(\next_ireg_3[14] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I10_G0N (.A(\un1_next_sum[10] )
        , .B(sum_10), .Y(N501));
    XNOR2 inf_abs1_a_2_I_28 (.A(sr_new[10]), .B(N_4), .Y(
        \inf_abs1_a_2[10] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I18_G0N (.A(
        \un1_next_sum_iv_1[18] ), .B(\un1_next_sum_iv_2[18] ), .C(
        sum_18), .Y(N525_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I338_un1_Y (.A(N846), .B(N877), 
        .Y(I338_un1_Y));
    DFN1E1C0 \p_adj[4]  (.D(\inf_abs1_5[4] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[4]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_2 (.A(
        ADD_22x22_fast_I144_un1_Y_0), .B(N425), .C(
        ADD_22x22_fast_I144_Y_1), .Y(ADD_22x22_fast_I144_Y_2));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I358_Y (.A(N878), .B(N743), .C(
        N877), .Y(N1073));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I7_G0N (.A(\i_adj[7]_net_1 ), 
        .B(\i_adj[9]_net_1 ), .Y(N287));
    XNOR2 inf_abs2_a_0_I_20 (.A(integral[13]), .B(N_20), .Y(
        \inf_abs2_a_0[7] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I424_Y_0 (.A(sum_6), .B(
        \un1_next_sum[6] ), .Y(ADD_40x40_fast_I424_Y_0));
    DFN1E1C0 \sumreg[17]  (.D(\next_sum[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_17));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I257_Y_1 (.A(N475), .B(N472), 
        .C(N661), .Y(ADD_40x40_fast_I257_Y_1));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I321_Y (.A(I321_un1_Y), .B(N815), 
        .Y(N1106));
    DFN1C0 \state[6]  (.D(\state[2]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[6]_net_1 ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I423_Y_0 (.A(
        \un1_next_sum_2[4] ), .B(\un1_next_sum_iv_0[5] ), .C(sum_5), 
        .Y(ADD_40x40_fast_I423_Y_0));
    AND3 inf_abs1_a_2_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[5] ), .Y(
        \DWACT_FINC_E[6] ));
    DFN1E1C0 \sumreg[35]  (.D(\next_sum[35] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[35]_net_1 ));
    MX2 \i_adj_RNO[13]  (.A(integral[19]), .B(\inf_abs2_a_0[13] ), .S(
        integral_1_0), .Y(\inf_abs2_5[13] ));
    DFN1E1C0 \sumreg[4]  (.D(\next_sum[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416), .Q(sum_4));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I87_un1_Y (.A(N358), .B(N266), 
        .Y(I87_un1_Y));
    XA1B \sumreg_RNO[38]  (.A(N1023), .B(ADD_40x40_fast_I456_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[38] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I160_Y (.A(N636), .B(N633), .C(
        N632), .Y(N713));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I232_Y (.A(N717), .B(N710), .C(
        N709), .Y(N791));
    NOR2 inf_abs2_a_0_I_6 (.A(integral[6]), .B(integral[7]), .Y(N_25));
    NOR3B inf_abs2_a_0_I_45 (.A(\DWACT_FINC_E[10] ), .B(
        \DWACT_FINC_E_0[6] ), .C(integral[21]), .Y(N_11_0));
    NOR3 inf_abs1_a_2_I_29 (.A(sr_new[7]), .B(sr_new[6]), .C(sr_new[8])
        , .Y(\DWACT_FINC_E_0[5] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I252_Y (.A(N737), .B(N730), .C(
        N729), .Y(N811));
    NOR3A \state_RNI0QFF[4]  (.A(integral[25]), .B(\state[5]_net_1 ), 
        .C(\state[4]_net_1 ), .Y(N_232));
    MX2 \p_adj_RNO[1]  (.A(sr_new[1]), .B(\inf_abs1_a_2[1] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[1] ));
    NOR3B \preg_RNI5OBI[11]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[11]_net_1 ), .Y(\un24_next_sum_m[11] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I382_un1_Y (.A(N878), .B(N743), 
        .C(N846), .Y(I382_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I53_Y (.A(N270), .B(N273), .Y(
        N358));
    AO1 next_ireg_3_0_ADD_22x22_fast_I30_Y (.A(N302), .B(N306), .C(
        N305), .Y(N335));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I124_un1_Y (.A(N377), .B(N369), 
        .C(N424), .Y(I124_un1_Y));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I330_un1_Y (.A(N770), .B(N754), 
        .C(N869), .Y(I330_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I237_Y (.A(N722), .B(N714), .Y(
        N796));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I12_G0N (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[12]_net_1 ), .Y(N302));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I11_G0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(N299));
    XA1 \ireg_RNI24NI[4]  (.A(integral_0_0), .B(\ireg[4]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[4] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I58_Y (.A(\sumreg[28]_net_1 ), 
        .B(\sumreg[29]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N608)
        );
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I257_Y (.A(
        ADD_40x40_fast_I257_Y_1), .B(N734), .Y(N816));
    OR2 \ireg_RNIEJPP1[6]  (.A(\un3_next_sum_m[6] ), .B(
        \un1_next_sum_iv_0[6] ), .Y(\un1_next_sum_iv_2[6] ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I35_Y (.A(\i_adj[10]_net_1 ), .B(
        \i_adj[12]_net_1 ), .C(N300), .Y(N340));
    NOR2B un1_sumreg_0_0_ADD_m8_i_a4_0_0 (.A(sum_0_d0), .B(sum_1_d0), 
        .Y(ADD_m8_i_a4_0_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I260_un1_Y (.A(N740), .B(N666), 
        .Y(I260_un1_Y));
    DFN1E1C0 \sumreg[7]  (.D(\next_sum[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416), .Q(sum_7));
    DFN1E1C0 \ireg[12]  (.D(\next_ireg_3[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[12]_net_1 ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I176_Y_0 (.A(\i_adj[16]_net_1 ), 
        .B(\i_adj[18]_net_1 ), .Y(ADD_22x22_fast_I176_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I126_Y (.A(N602), .B(N598), .Y(
        N679));
    NOR2A inf_abs2_a_0_I_11 (.A(\DWACT_FINC_E_0[0] ), .B(integral[9]), 
        .Y(N_23));
    OR2 \state_RNIQSHS[5]  (.A(next_sum_0_sqmuxa_1), .B(
        next_sum_0_sqmuxa_2), .Y(\un1_next_sum_2[4] ));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I166_Y (.A(\i_adj[8]_net_1 ), .B(
        \i_adj[6]_net_1 ), .C(N528), .Y(\next_ireg_3[12] ));
    NOR2B \preg_RNICVBI_0[18]  (.A(\preg[18]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[18] ));
    OA1A un1_sumreg_0_0_ADD_40x40_fast_I67_Y (.A(
        \un1_next_sum_0_iv[25] ), .B(\sumreg[25]_net_1 ), .C(N544), .Y(
        N617));
    AO1 next_ireg_3_0_ADD_22x22_fast_I38_Y (.A(N290), .B(N294), .C(
        N293), .Y(N343));
    XNOR2 inf_abs2_a_0_I_46 (.A(integral[22]), .B(N_11_0), .Y(
        \inf_abs2_a_0[16] ));
    XOR2 inf_abs1_a_2_I_5 (.A(sr_new[0]), .B(sr_new[1]), .Y(
        \inf_abs1_a_2[1] ));
    XNOR2 inf_abs1_a_2_I_23 (.A(sr_new[8]), .B(N_6_0), .Y(
        \inf_abs1_a_2[8] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I310_Y (.A(N813), .B(N798), .C(
        N797), .Y(N881));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I169_Y (.A(N645), .B(N641), .Y(
        N722));
    DFN1C0 \state[2]  (.D(\state[1]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[2]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I245_Y (.A(N730), .B(N722), .Y(
        N804));
    DFN1E1C0 \i_adj[15]  (.D(\inf_abs2_5[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[15]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I41_Y (.A(N291), .B(N288), .Y(
        N346));
    DFN1E1C0 \i_adj[20]  (.D(\inf_abs2_5[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[20]_net_1 ));
    XNOR2 inf_abs2_a_0_I_37 (.A(integral[19]), .B(N_14), .Y(
        \inf_abs2_a_0[13] ));
    MX2 \i_adj_RNO[12]  (.A(integral[18]), .B(\inf_abs2_a_0[12] ), .S(
        integral_1_0), .Y(\inf_abs2_5[12] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I53_Y (.A(\sumreg[32]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N603)
        );
    OR2 next_ireg_3_0_ADD_22x22_fast_I86_Y (.A(I86_un1_Y), .B(N355), 
        .Y(N394));
    AX1D next_ireg_3_0_ADD_22x22_fast_I170_Y (.A(N422), .B(I132_un1_Y), 
        .C(ADD_22x22_fast_I170_Y_0), .Y(\next_ireg_3[16] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_1 (.A(N369), .B(N376), .C(
        ADD_22x22_fast_I144_Y_0), .Y(ADD_22x22_fast_I144_Y_1));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I4_P0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[4] ), .C(sum_4), .Y(N484));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I213_Y (.A(N690), .B(N698), .Y(
        N772));
    DFN1E1C0 \p_adj[10]  (.D(\inf_abs1_5[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[10]_net_1 ));
    DFN1E1C0 \p_adj[5]  (.D(\inf_abs1_5[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[5]_net_1 ));
    NOR3B \preg_RNI6PBI[12]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[12]_net_1 ), .Y(\un24_next_sum_m[12] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I164_Y (.A(N640), .B(N637), .C(
        N636), .Y(N717));
    DFN1E1C0 \sumreg[36]  (.D(\next_sum[36] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[36]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I56_Y (.A(\sumreg[29]_net_1 ), 
        .B(\sumreg[30]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N606)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I172_Y (.A(N648), .B(N645), .C(
        N644), .Y(N725));
    NOR2B \p_adj_RNO[12]  (.A(\inf_abs1_a_2[12] ), .B(sr_new[12]), .Y(
        \inf_abs1_5[12] ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I126_un1_Y (.A(N386), .B(
        I112_un1_Y), .C(ADD_22x22_fast_I126_un1_Y_0), .Y(I126_un1_Y));
    NOR3B \ireg_RNI8P101[18]  (.A(integral_0_0), .B(\state[3]_net_1 ), 
        .C(\ireg[18]_net_1 ), .Y(\un3_next_sum_m[18] ));
    DFN1E1C0 \p_adj[0]  (.D(\inf_abs1_5[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[0]_net_1 ));
    AND3 inf_abs2_a_0_I_51 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[28] ));
    OR2 \preg_RNINV3M3[10]  (.A(\un1_next_sum_iv_2[10] ), .B(
        \un1_next_sum_iv_1[10] ), .Y(\un1_next_sum[10] ));
    DFN1E1C0 \sumreg[9]  (.D(\next_sum[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416), .Q(sum_9));
    NOR3B \preg_RNICLDK[9]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[9]_net_1 ), .Y(\un24_next_sum_m[9] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I181_Y (.A(N657), .B(N653), .Y(
        N734));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I216_Y (.A(N701), .B(N694), .C(
        N693), .Y(N775));
    OA1 un1_sumreg_0_0_ADD_m8_i_a4 (.A(N_232), .B(ADD_m8_i_o4_1), .C(
        next_sum_0_sqmuxa), .Y(ADD_m8_i_a4));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I4_G0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[4] ), .C(sum_4), .Y(N483));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I317_Y (.A(N808), .B(N823), .C(
        N807), .Y(N1094));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I129_Y (.A(N601), .B(N605), .Y(
        N682));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I50_Y (.A(N272), .B(
        \i_adj[3]_net_1 ), .C(\i_adj[5]_net_1 ), .Y(N355));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I144_un1_Y_0 (.A(N377), .B(N369)
        , .C(N266), .Y(ADD_22x22_fast_I144_un1_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I34_Y (.A(N296), .B(N300), .C(
        N299), .Y(N339));
    DFN1E1C0 \sumreg[31]  (.D(\next_sum[31] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[31]_net_1 ));
    DFN1E1C0 \sumreg[2]  (.D(\next_sum[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416), .Q(sum_2_d0));
    DFN1E1C0 \i_adj[7]  (.D(\inf_abs2_5[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[7]_net_1 ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I383_Y (.A(
        ADD_40x40_fast_I383_Y_1), .B(I383_un1_Y), .C(I340_un1_Y), .Y(
        N1031));
    MX2 \i_adj_RNO[8]  (.A(integral[14]), .B(\inf_abs2_a_0[8] ), .S(
        integral[25]), .Y(\inf_abs2_5[8] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I9_P0N (.A(
        \un1_next_sum_iv_1[9] ), .B(\un1_next_sum_iv_2[9] ), .C(sum_9), 
        .Y(N499));
    OR2 \ireg_RNICMRG3[15]  (.A(\un1_next_sum_iv_2[15] ), .B(
        \un1_next_sum_iv_1[15] ), .Y(\un1_next_sum[15] ));
    NOR3A inf_abs2_a_0_I_27 (.A(\DWACT_FINC_E_0[4] ), .B(integral[14]), 
        .C(integral[15]), .Y(N_17));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I105_Y (.A(sum_6), .B(
        \un1_next_sum[6] ), .C(N487), .Y(N655));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I10_G0N (.A(\i_adj[12]_net_1 ), 
        .B(\i_adj[10]_net_1 ), .Y(N296));
    AO1 next_ireg_3_0_ADD_22x22_fast_I108_Y (.A(N390), .B(N383), .C(
        N382), .Y(N422));
    MX2 \p_adj_RNO[3]  (.A(sr_new[3]), .B(\inf_abs1_a_2[3] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[3] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I435_Y_0 (.A(sum_17), .B(
        \un1_next_sum[17] ), .Y(ADD_40x40_fast_I435_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I146_Y (.A(N622), .B(N619), .C(
        N618), .Y(N699));
    NOR3B \preg_RNI4NBI[10]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[10]_net_1 ), .Y(\un24_next_sum_m[10] ));
    OR2 \preg_RNI3C361[10]  (.A(next_sum_0_sqmuxa_1), .B(
        \un24_next_sum_m[10] ), .Y(\un1_next_sum_iv_0[10] ));
    AND3 inf_abs2_a_0_I_48 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[11] ), .Y(N_10_0));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I197_Y_0 (.A(\sumreg[37]_net_1 )
        , .B(\sumreg[36]_net_1 ), .C(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I197_Y_0));
    DFN1E1C0 \preg[16]  (.D(\p_adj[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[16]_net_1 ));
    NOR3 \state_RNI8K6L[6]  (.A(sum_rdy), .B(\state[6]_net_1 ), .C(
        \state[1]_net_1 ), .Y(N_416));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I135_Y (.A(N607), .B(N611), .Y(
        N688));
    DFN1E1C0 \preg[17]  (.D(\p_adj[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[17]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I9_G0N (.A(\i_adj[11]_net_1 ), 
        .B(\i_adj[9]_net_1 ), .Y(N293));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I155_Y (.A(N627), .B(N631), .Y(
        N708));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I122_un1_Y (.A(N407), .B(N422), 
        .Y(I122_un1_Y));
    NOR3B \preg_RNIBUBI[17]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[17]_net_1 ), .Y(\un24_next_sum_m[17] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I5_P0N (.A(\i_adj[7]_net_1 ), .B(
        \i_adj[5]_net_1 ), .Y(N282));
    DFN1E1C0 \i_adj[8]  (.D(\inf_abs2_5[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[8]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I94_Y (.A(N501), .B(N505), .C(
        N504_0), .Y(N644));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I73_Y (.A(N342), .B(N346), .Y(
        N381));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I174_Y (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .C(N504), .Y(\next_ireg_3[20] ));
    DFN1E1C0 \i_adj[17]  (.D(\inf_abs2_5[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[17]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I214_un1_Y (.A(N699), .B(N692), 
        .Y(I214_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I140_Y (.A(N616), .B(N613), .C(
        N612), .Y(N693));
    MX2 \i_adj_RNO[3]  (.A(integral[9]), .B(\inf_abs2_a_0[3] ), .S(
        integral_1_0), .Y(\inf_abs2_5[3] ));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I74_Y (.A(N531_0), .B(sum_21), 
        .C(\un1_next_sum[21] ), .Y(N624));
    XNOR2 inf_abs2_a_0_I_49 (.A(integral[23]), .B(N_10_0), .Y(
        \inf_abs2_a_0[17] ));
    XNOR2 inf_abs2_a_0_I_12 (.A(integral[10]), .B(N_23), .Y(
        \inf_abs2_a_0[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I319_Y (.A(N812), .B(N745), .C(
        N811), .Y(N1100));
    XA1B \sumreg_RNO[18]  (.A(N1076), .B(ADD_40x40_fast_I436_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[18] ));
    NOR3B \ireg_RNIG8DP[11]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[11]_net_1 ), .Y(\un3_next_sum_m[11] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I306_Y (.A(N809), .B(N794), .C(
        N793), .Y(N877));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I224_Y (.A(N709), .B(N702), .C(
        N701), .Y(N783));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I209_Y (.A(N686), .B(N694), .Y(
        N768));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I383_Y_0 (.A(N681), .B(N689), .Y(
        ADD_40x40_fast_I383_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I17_G0N (.A(\un1_next_sum[17] )
        , .B(sum_17), .Y(N522));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I356_Y (.A(N874), .B(N821), .C(
        N873), .Y(N1067));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I239_Y (.A(N724), .B(N716), .Y(
        N798));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I259_Y (.A(N738), .B(N745), .C(
        N737), .Y(N819));
    NOR2B \i_adj_RNO[21]  (.A(\inf_abs2_a_0[21] ), .B(integral[25]), 
        .Y(\inf_abs2_5[21] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I116_un1_Y (.A(N472), .B(
        \un1_next_sum[0] ), .Y(I116_un1_Y));
    DFN1E1C0 \sumreg[6]  (.D(\next_sum[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416), .Q(sum_6));
    DFN1E1C0 \sumreg[0]  (.D(\next_sum[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416), .Q(sum_0_d0));
    DFN1E1C0 \preg[15]  (.D(\p_adj[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[15]_net_1 ));
    DFN1E1C0 \i_adj[10]  (.D(\inf_abs2_5[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[10]_net_1 ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I452_Y_0 (.A(
        \sumreg[34]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I452_Y_0));
    DFN1E1C0 \ireg[24]  (.D(\next_ireg_3[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[24]_net_1 ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I351_un1_Y (.A(N780), .B(N796), 
        .C(N1100), .Y(I351_un1_Y));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I347_un1_Y (.A(N772), .B(N788), 
        .C(N1088), .Y(I347_un1_Y));
    XNOR2 inf_abs2_a_0_I_43 (.A(integral[21]), .B(N_12_0), .Y(
        \inf_abs2_a_0[15] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I69_Y (.A(N338), .B(N342), .Y(
        N377));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I385_Y (.A(I385_un1_Y), .B(
        ADD_40x40_fast_I385_Y_1), .C(I344_un1_Y), .Y(N1035));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I149_Y (.A(N621), .B(N625), .Y(
        N702));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I67_Y (.A(N336), .B(N340), .Y(
        N375));
    OR2 next_ireg_3_0_ADD_22x22_fast_I54_Y (.A(I87_un1_Y), .B(N269), 
        .Y(N359));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I378_Y_2 (.A(N594), .B(
        ADD_40x40_fast_I378_Y_0), .C(N679), .Y(ADD_40x40_fast_I378_Y_2)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I360_Y (.A(N882), .B(N666), .C(
        N881), .Y(N1079));
    MX2 \p_adj_RNO[0]  (.A(sr_new[0]), .B(sr_new[0]), .S(sr_new_0_0), 
        .Y(\inf_abs1_5[0] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I384_Y_0 (.A(N691), .B(N684), .C(
        N683), .Y(ADD_40x40_fast_I384_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I182_Y (.A(N658), .B(N655), .C(
        N654), .Y(N735));
    AND3 inf_abs2_a_0_I_52 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[12] ), .Y(N_9_0));
    NOR3A inf_abs2_a_0_I_31 (.A(\DWACT_FINC_E_0[6] ), .B(integral[15]), 
        .C(integral[16]), .Y(N_16));
    NOR3B \ireg_RNI8EKH[8]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[8]_net_1 ), .Y(\un3_next_sum_m[8] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I163_Y (.A(N639), .B(N635), .Y(
        N716));
    AO1 next_ireg_3_0_ADD_22x22_fast_I110_Y (.A(N392), .B(N385), .C(
        N384), .Y(N424));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I197_Y (.A(N597), .B(
        ADD_40x40_fast_I197_Y_0), .C(N682), .Y(N756));
    DFN1E1C0 \i_adj[18]  (.D(\inf_abs2_5[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[18]_net_1 ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I91_Y (.A(sum_12), .B(
        \un1_next_sum[12] ), .C(N511), .Y(N641));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I93_Y (.A(N367), .B(N375), .Y(
        N407));
    OR2 \ireg_RNIB70M1[21]  (.A(\un1_next_sum_iv_0[21] ), .B(
        \un1_next_sum_2[4] ), .Y(\un1_next_sum[21] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I144_Y (.A(N620), .B(N617), .C(
        N616), .Y(N697));
    MX2 \i_adj_RNO[16]  (.A(integral[22]), .B(\inf_abs2_a_0[16] ), .S(
        integral_1_0), .Y(\inf_abs2_5[16] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I71_Y (.A(N541), .B(N538), .Y(
        N621));
    NOR3B \ireg_RNI57NI[7]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[7]_net_1 ), .C(integral_0_0), .Y(\ireg_m[7] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I95_Y (.A(sum_10), .B(
        \un1_next_sum[10] ), .C(N505), .Y(N645));
    OR2 next_ireg_3_0_ADD_22x22_fast_I13_P0N (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[13]_net_1 ), .Y(N306));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I161_Y (.A(\i_adj[3]_net_1 ), .B(
        \i_adj[1]_net_1 ), .C(N266), .Y(\next_ireg_3[7] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I70_Y (.A(N343), .B(N340), .C(
        N339), .Y(N378));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I75_Y (.A(sum_21), .B(
        \un1_next_sum[21] ), .C(N532), .Y(N625));
    OR3 \preg_RNIOPGV1[13]  (.A(\un24_next_sum_m[13] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[13] ), .Y(
        \un1_next_sum_iv_2[13] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I168_Y (.A(N644), .B(N641), .C(
        N640), .Y(N721));
    MX2 \p_adj_RNO[6]  (.A(sr_new[6]), .B(\inf_abs1_a_2[6] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[6] ));
    AO1 \ireg_RNI1HMA1[16]  (.A(\ireg[16]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[16] ), .Y(
        \un1_next_sum_iv_1[16] ));
    MX2 \i_adj_RNO[1]  (.A(integral[7]), .B(\inf_abs2_a_0[1] ), .S(
        integral_1_0), .Y(\inf_abs2_5[1] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I75_Y (.A(N348), .B(N344), .Y(
        N383));
    GND GND_i (.Y(GND));
    NOR2A \state_RNIR7Q8_0[5]  (.A(\state[5]_net_1 ), .B(sr_new[12]), 
        .Y(next_sum_1_sqmuxa_2));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I143_Y_0 (.A(\i_adj[17]_net_1 ), 
        .B(\i_adj[19]_net_1 ), .C(N314), .Y(ADD_22x22_fast_I143_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I244_Y (.A(N729), .B(N722), .C(
        N721), .Y(N803));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I314_Y (.A(N802), .B(N817), .C(
        N801), .Y(N1085));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I320_Y (.A(N814), .B(N666), .C(
        N813), .Y(N1103));
    NOR3B \ireg_RNI3N741[12]  (.A(\state[3]_net_1 ), .B(
        \ireg[12]_net_1 ), .C(integral_1_0), .Y(\ireg_m[12] ));
    MX2 \p_adj_RNO[5]  (.A(sr_new[5]), .B(\inf_abs1_a_2[5] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[5] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I378_Y_3 (.A(N754), .B(N769), .C(
        ADD_40x40_fast_I378_Y_2), .Y(ADD_40x40_fast_I378_Y_3));
    DFN1C0 \state[5]  (.D(\state[4]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[5]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I78_Y (.A(N351), .B(N348), .C(
        N347), .Y(N386));
    NOR2 inf_abs2_a_0_I_21 (.A(integral[13]), .B(integral[12]), .Y(
        \DWACT_FINC_E[3] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I418_Y_0 (.A(sum_0_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I418_Y_0));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I87_Y (.A(sum_15), .B(
        \un1_next_sum[15] ), .C(N514), .Y(N637));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I384_Y_2 (.A(
        ADD_40x40_fast_I384_Y_0), .B(I278_un1_Y), .C(I384_un1_Y), .Y(
        ADD_40x40_fast_I384_Y_2));
    OA1 next_ireg_3_0_ADD_22x22_fast_I29_Y (.A(\i_adj[16]_net_1 ), .B(
        \i_adj[14]_net_1 ), .C(N306), .Y(N334));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I22_P0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[22] ), .C(sum_22), .Y(N538));
    NOR3A inf_abs1_a_2_I_31 (.A(\DWACT_FINC_E[6] ), .B(sr_new[9]), .C(
        sr_new[10]), .Y(N_3));
    OA1 next_ireg_3_0_ADD_22x22_fast_I27_Y (.A(\i_adj[16]_net_1 ), .B(
        \i_adj[14]_net_1 ), .C(N312), .Y(N332));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I223_Y (.A(N700), .B(N708), .Y(
        N782));
    DFN1E1C0 \ireg[6]  (.D(\next_ireg_3[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[6]_net_1 ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I334_un1_Y (.A(N774), .B(N758), 
        .C(N873), .Y(I334_un1_Y));
    OR3 \preg_RNID7562[15]  (.A(\un24_next_sum_m[15] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[15] ), .Y(
        \un1_next_sum_iv_2[15] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I23_G0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[23] ), .C(sum_23), .Y(N540));
    DFN1E1C0 \preg[6]  (.D(\p_adj[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[6]_net_1 ));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I36_Y (.A(N293), .B(
        \i_adj[10]_net_1 ), .C(\i_adj[12]_net_1 ), .Y(N341));
    NOR2 inf_abs1_a_2_I_6 (.A(sr_new[0]), .B(sr_new[1]), .Y(N_12));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I1_G0N (.A(\i_adj[1]_net_1 ), 
        .B(\i_adj[3]_net_1 ), .Y(N269));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I318_Y (.A(I318_un1_Y), .B(N809), 
        .Y(N1097));
    AO1 next_ireg_3_0_ADD_22x22_fast_I114_Y (.A(N391), .B(N359), .C(
        N390), .Y(N528));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I64_Y (.A(I64_un1_Y), .B(N549), 
        .Y(N614));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I457_Y_0 (.A(sum_39), .B(
        \un1_next_sum_1_iv[26] ), .Y(ADD_40x40_fast_I457_Y_0));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I186_un1_Y (.A(N484), .B(N481), 
        .C(N662), .Y(I186_un1_Y));
    XA1B \sumreg_RNO[34]  (.A(N1031), .B(ADD_40x40_fast_I452_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[34] ));
    XA1 \ireg_RNIG9EP[20]  (.A(integral_0_0), .B(\ireg[20]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[20] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I81_Y (.A(N354), .B(N350), .Y(
        N389));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I128_Y (.A(N604), .B(N600), .Y(
        N681));
    NOR3B \preg_RNIATBI[16]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[16]_net_1 ), .Y(\un24_next_sum_m[16] ));
    DFN1E1C0 \sumreg[29]  (.D(\next_sum[29] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[29]_net_1 ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I99_Y (.A(sum_8), .B(
        \un1_next_sum[8] ), .C(N499), .Y(N649));
    OR2 \ireg_RNIN87A3[14]  (.A(\un1_next_sum_iv_2[14] ), .B(
        \un1_next_sum_iv_1[14] ), .Y(\un1_next_sum[14] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I169_Y_0 (.A(\i_adj[9]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(ADD_22x22_fast_I169_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I226_Y (.A(N711), .B(N704), .C(
        N703), .Y(N785));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I442_Y_0 (.A(
        \un1_next_sum_2[4] ), .B(\un1_next_sum_iv_0[24] ), .C(
        \sumreg[24]_net_1 ), .Y(ADD_40x40_fast_I442_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I212_Y (.A(N697), .B(N690), .C(
        N689), .Y(N771));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I79_Y (.A(sum_19), .B(
        \un1_next_sum[19] ), .C(N526), .Y(N629));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I167_Y (.A(N639), .B(N643), .Y(
        N720));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I164_Y_0 (.A(\i_adj[4]_net_1 ), 
        .B(\i_adj[6]_net_1 ), .Y(ADD_22x22_fast_I164_Y_0));
    NOR3 inf_abs1_a_2_I_10 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2])
        , .Y(\DWACT_FINC_E[0] ));
    DFN1C0 \state_0[3]  (.D(\state[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_0[3]_net_1 ));
    DFN1E1C0 \ireg[21]  (.D(\next_ireg_3[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[21]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I281_Y (.A(N768), .B(N784), .Y(
        N852));
    AO1 \preg_RNI3R241[9]  (.A(\preg[9]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[9] ), .Y(
        \un1_next_sum_iv_1[9] ));
    XNOR2 inf_abs2_a_0_I_32 (.A(integral[17]), .B(N_16), .Y(
        \inf_abs2_a_0[11] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I430_Y_0 (.A(sum_12), .B(
        \un1_next_sum[12] ), .Y(ADD_40x40_fast_I430_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I217_Y (.A(N702), .B(N694), .Y(
        N776));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I378_un1_Y (.A(N770), .B(N754), 
        .C(ADD_40x40_fast_I378_un1_Y_0), .Y(I378_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I275_Y (.A(N762), .B(N778), .Y(
        N846));
    XA1B \sumreg_RNO[27]  (.A(N1049), .B(ADD_40x40_fast_I445_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[27] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I74_Y (.A(N347), .B(N344), .C(
        N343), .Y(N382));
    DFN1E1C0 \sumreg[19]  (.D(\next_sum[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_19));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I422_Y_0 (.A(
        \un1_next_sum_2[4] ), .B(\un1_next_sum_iv_0[4] ), .C(sum_4), 
        .Y(ADD_40x40_fast_I422_Y_0));
    DFN1E1C0 \sumreg[8]  (.D(\next_sum[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416), .Q(sum_8));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I349_un1_Y (.A(N776), .B(N792), 
        .C(N1094), .Y(I349_un1_Y));
    DFN1E1C0 \sumreg[28]  (.D(\next_sum[28] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[28]_net_1 ));
    AO1A \state_RNIQSHS[4]  (.A(derivative_0), .B(\state[4]_net_1 ), 
        .C(next_sum_1_sqmuxa_2), .Y(\un1_next_sum_0_iv_0[25] ));
    XA1B \sumreg_RNO[0]  (.A(N_228), .B(ADD_40x40_fast_I418_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[0] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I451_Y_0 (.A(
        \sumreg[33]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I451_Y_0));
    XA1 \ireg_RNIJCEP[23]  (.A(integral_0_0), .B(\ireg[23]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[23] ));
    OR3 \preg_RNIGLPP1[7]  (.A(\un24_next_sum_m[7] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[7] ), .Y(
        \un1_next_sum_iv_2[7] ));
    AO1 \preg_RNIVM241[7]  (.A(\preg[7]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[7] ), .Y(
        \un1_next_sum_iv_1[7] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_1_0 (.A(
        ADD_22x22_fast_I142_Y_0_a3_0), .B(N330), .Y(
        ADD_22x22_fast_I142_Y_0_a3_1));
    DFN1C0 \state_2[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_2[2]_net_1 ));
    DFN1E1C0 \sumreg[18]  (.D(\next_sum[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_18));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I380_Y_1 (.A(N598), .B(N594), .C(
        N683), .Y(ADD_40x40_fast_I380_Y_1));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I61_Y (.A(\sumreg[28]_net_1 ), 
        .B(\sumreg[27]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N611)
        );
    OR2 \state_RNI9CV41_0[4]  (.A(\un1_next_sum_0_iv_0[25] ), .B(
        next_sum_1_sqmuxa), .Y(\un1_next_sum_1_iv[26] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I6_G0N (.A(\i_adj[8]_net_1 ), 
        .B(\i_adj[6]_net_1 ), .Y(N284));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I162_Y (.A(
        ADD_22x22_fast_I162_Y_0), .B(N359), .Y(\next_ireg_3[8] ));
    NOR2B \ireg_RNINKBO[25]  (.A(\ireg[25]_net_1 ), .B(
        next_sum_0_sqmuxa), .Y(\ireg_m[25] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I243_Y (.A(N720), .B(N728), .Y(
        N802));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I127_Y (.A(N599), .B(N603), .Y(
        N680));
    DFN1E1C0 \p_adj[3]  (.D(\inf_abs1_5[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[3]_net_1 ));
    DFN1E1C0 \ireg[10]  (.D(\next_ireg_3[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[10]_net_1 ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I49_Y (.A(\i_adj[3]_net_1 ), .B(
        \i_adj[5]_net_1 ), .C(N279), .Y(N354));
    OA1A un1_sumreg_0_0_ADD_40x40_fast_I65_Y (.A(
        \un1_next_sum_0_iv[25] ), .B(\sumreg[25]_net_1 ), .C(N550), .Y(
        N615));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I47_Y (.A(N282), .B(N279), .Y(
        N352));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I101_Y (.A(sum_8), .B(
        \un1_next_sum[8] ), .C(N493), .Y(N651));
    AND3 inf_abs2_a_0_I_22 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_19));
    DFN1E1C0 \sumreg[1]  (.D(\next_sum[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416), .Q(sum_1_d0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I449_Y_0 (.A(
        \sumreg[31]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I449_Y_0));
    XA1B \sumreg_RNO[20]  (.A(N1070), .B(ADD_40x40_fast_I438_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[20] ));
    DFN1E1C0 \sumreg_0[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(sum_0_0));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I47_Y (.A(\sumreg[35]_net_1 ), 
        .B(\sumreg[34]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N597)
        );
    XNOR2 inf_abs1_a_2_I_32 (.A(sr_new[11]), .B(N_3), .Y(
        \inf_abs1_a_2[11] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I187_Y_0 (.A(\un1_next_sum[0] ), 
        .B(sum_2_d0), .C(N475), .Y(ADD_40x40_fast_I187_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I148_Y (.A(N624), .B(N621), .C(
        N620), .Y(N701));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I165_Y (.A(
        ADD_22x22_fast_I165_Y_0), .B(N531), .Y(\next_ireg_3[11] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I13_G0N (.A(\un1_next_sum[13] )
        , .B(sum_13), .Y(N510_0));
    XA1B \sumreg_RNO[21]  (.A(N1067), .B(ADD_40x40_fast_I439_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[21] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_3_0 (.A(N338), .B(
        N334), .Y(ADD_22x22_fast_I142_Y_0_a3_3_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I131_Y (.A(N603), .B(N607), .Y(
        N684));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I86_un1_Y (.A(N356), .B(N359), 
        .Y(I86_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I303_Y (.A(N806), .B(N790), .Y(
        N874));
    XNOR2 inf_abs1_a_2_I_20 (.A(sr_new[7]), .B(N_7_1), .Y(
        \inf_abs1_a_2[7] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I438_Y_0 (.A(
        \un1_next_sum_2[4] ), .B(\un1_next_sum_iv_0[20] ), .C(sum_20), 
        .Y(ADD_40x40_fast_I438_Y_0));
    DFN1E1C0 \sumreg[25]  (.D(\next_sum[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[25]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I246_Y (.A(N731), .B(N724), .C(
        N723), .Y(N805));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I151_Y (.A(N623), .B(N627), .Y(
        N704));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I176_Y (.A(N652), .B(N649), .C(
        N648), .Y(N729));
    OR2 \state_RNI9CV41[3]  (.A(\un1_next_sum_2[4] ), .B(
        next_sum_0_sqmuxa), .Y(\un1_next_sum[0] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I347_Y (.A(
        ADD_40x40_fast_I347_Y_0), .B(I347_un1_Y), .Y(N1040));
    DFN1E1C0 \ireg[23]  (.D(\next_ireg_3[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[23]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I106_un1_Y (.A(N381), .B(N388), 
        .Y(I106_un1_Y));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I429_Y_0 (.A(sum_11), .B(
        \un1_next_sum[11] ), .Y(ADD_40x40_fast_I429_Y_0));
    OR3 un1_sumreg_0_0_ADD_m8_i (.A(ADD_m8_i_a4_0), .B(
        \un1_next_sum_2[4] ), .C(ADD_m8_i_a4), .Y(N743));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I9_G0N (.A(
        \un1_next_sum_iv_1[9] ), .B(\un1_next_sum_iv_2[9] ), .C(sum_9), 
        .Y(N498));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I447_Y_0 (.A(
        \sumreg[29]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I447_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I353_Y (.A(
        ADD_40x40_fast_I353_un1_Y_0), .B(N1106), .C(
        ADD_40x40_fast_I353_Y_0), .Y(N1058));
    AO1 \preg_RNI9GJM1[12]  (.A(\preg[12]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[12] ), .Y(
        \un1_next_sum_iv_1[12] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I379_Y_4 (.A(I268_un1_Y), .B(
        ADD_40x40_fast_I379_Y_2), .C(I332_un1_Y), .Y(
        ADD_40x40_fast_I379_Y_4));
    AND3 inf_abs2_a_0_I_60 (.A(integral_i[24]), .B(integral_i[25]), .C(
        integral_i[25]), .Y(\DWACT_FINC_E[15] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I170_Y (.A(N646), .B(N643), .C(
        N642), .Y(N723));
    DFN1E1C0 \sumreg[15]  (.D(\next_sum[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_15));
    DFN1E1C0 \ireg[5]  (.D(\i_adj[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[5]_net_1 ));
    DFN1E1C0 \ireg[25]  (.D(\next_ireg_3[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[25]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0 (.A(
        ADD_22x22_fast_I142_Y_0_a3_1), .B(N_11), .C(
        ADD_22x22_fast_I142_Y_0_1), .Y(N492));
    AO1 \preg_RNI7EJM1[11]  (.A(\preg[11]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[11] ), .Y(
        \un1_next_sum_iv_1[11] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I353_Y_0 (.A(N799), .B(N784), .C(
        N783), .Y(ADD_40x40_fast_I353_Y_0));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I5_G0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[5] ), .C(sum_5), .Y(N486));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I427_Y_0 (.A(
        \un1_next_sum_iv_1[9] ), .B(\un1_next_sum_iv_2[9] ), .C(sum_9), 
        .Y(ADD_40x40_fast_I427_Y_0));
    DFN1E1C0 \p_adj[9]  (.D(\inf_abs1_5[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[9]_net_1 ));
    XNOR2 inf_abs1_a_2_I_17 (.A(sr_new[6]), .B(N_8_0), .Y(
        \inf_abs1_a_2[6] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I163_Y (.A(
        ADD_22x22_fast_I163_Y_0), .B(N396), .Y(\next_ireg_3[9] ));
    MX2 \i_adj_RNO[14]  (.A(integral[20]), .B(\inf_abs2_a_0[14] ), .S(
        integral_1_0), .Y(\inf_abs2_5[14] ));
    NOR3B \ireg_RNI6N101[16]  (.A(integral_0_0), .B(\state[3]_net_1 ), 
        .C(\ireg[16]_net_1 ), .Y(\un3_next_sum_m[16] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I69_Y (.A(N541), .B(N544), .Y(
        N619));
    XA1B \sumreg_RNO[14]  (.A(N1088), .B(ADD_40x40_fast_I432_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[14] ));
    NOR2A \state_RNIFFD8_0[3]  (.A(\state[3]_net_1 ), .B(integral[25]), 
        .Y(next_sum_1_sqmuxa));
    XA1B \sumreg_RNO[35]  (.A(N1029), .B(ADD_40x40_fast_I453_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[35] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I349_Y (.A(I288_un1_Y), .B(N775), 
        .C(I349_un1_Y), .Y(N1046));
    DFN1C0 \state[4]  (.D(\state[3]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[4]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I147_Y (.A(N619), .B(N623), .Y(
        N700));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I8_G0N (.A(\i_adj[8]_net_1 ), 
        .B(\i_adj[10]_net_1 ), .Y(N290));
    AO13 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_0 (.A(\i_adj[20]_net_1 )
        , .B(\i_adj[18]_net_1 ), .C(N_7), .Y(ADD_22x22_fast_I142_Y_0_0)
        );
    AO1 \preg_RNITK241[6]  (.A(\preg[6]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[6] ), .Y(
        \un1_next_sum_iv_1[6] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I9_P0N (.A(\i_adj[11]_net_1 ), .B(
        \i_adj[9]_net_1 ), .Y(N294));
    NOR2A \ireg_RNINKBO_0[25]  (.A(next_sum_1_sqmuxa), .B(
        \ireg[25]_net_1 ), .Y(\un3_next_sum_m[25] ));
    DFN1E1C0 \sumreg[26]  (.D(\next_sum[26] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[26]_net_1 ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I441_Y_0 (.A(
        \un1_next_sum_2[4] ), .B(\un1_next_sum_iv_0[23] ), .C(sum_23), 
        .Y(ADD_40x40_fast_I441_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I179_Y (.A(N651), .B(N655), .Y(
        N732));
    XA1B \sumreg_RNO[7]  (.A(N817), .B(ADD_40x40_fast_I425_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[7] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I11_P0N (.A(\un1_next_sum[11] ), 
        .B(sum_11), .Y(N505));
    OR2 \preg_RNIAJ361[17]  (.A(next_sum_0_sqmuxa_1), .B(
        \un24_next_sum_m[17] ), .Y(\un1_next_sum_iv_0[17] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I128_Y_0 (.A(N382), .B(N375), .C(
        N374), .Y(ADD_22x22_fast_I128_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I90_Y (.A(N507_0), .B(N511), .C(
        N510_0), .Y(N640));
    DFN1E1C0 \ireg[17]  (.D(\next_ireg_3[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[17]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I316_Y (.A(N806), .B(N821), .C(
        N805), .Y(N1091));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I305_Y (.A(N808), .B(N792), .Y(
        N876));
    OR2 \preg_RNIJGST2[8]  (.A(\un1_next_sum_iv_2[8] ), .B(
        \un1_next_sum_iv_1[8] ), .Y(\un1_next_sum[8] ));
    NOR2B \state_RNIVKNJ[4]  (.A(\state[4]_net_1 ), .B(derivative_0), 
        .Y(next_sum_0_sqmuxa_1));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I381_Y (.A(
        ADD_40x40_fast_I381_Y_2), .B(I381_un1_Y), .C(I336_un1_Y), .Y(
        N1027));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I219_Y (.A(N619), .B(N615), .C(
        N704), .Y(N778));
    XA1 \ireg_RNIIBEP[22]  (.A(integral_0_0), .B(\ireg[22]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[22] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I102_Y (.A(N489), .B(N493), .C(
        N492_0), .Y(N652));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I70_Y (.A(N537), .B(N541), .C(
        N540), .Y(N620));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I21_G0N (.A(\un1_next_sum[21] )
        , .B(sum_21), .Y(N534));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I195_Y (.A(N595), .B(
        ADD_40x40_fast_I195_Y_0), .C(N680), .Y(N754));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I421_Y_0 (.A(sum_3), .B(N743), 
        .Y(ADD_40x40_fast_I421_Y_0));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I318_un1_Y (.A(N728), .B(N736), 
        .C(N743), .Y(I318_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I174_Y (.A(N650), .B(N647), .C(
        N646), .Y(N727));
    DFN1E1C0 \sumreg[16]  (.D(\next_sum[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_16));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I16_G0N (.A(\i_adj[18]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .Y(N314));
    XNOR2 inf_abs2_a_0_I_14 (.A(integral[11]), .B(N_22), .Y(
        \inf_abs2_a_0[5] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I355_Y (.A(N872), .B(N819), .C(
        N871), .Y(N1064));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I132_Y (.A(N608), .B(N604), .Y(
        N685));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I2_G0N (.A(\i_adj[2]_net_1 ), 
        .B(\i_adj[4]_net_1 ), .Y(N272));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I152_Y (.A(N628), .B(N625), .C(
        N624), .Y(N705));
    MX2 \p_adj_RNO[8]  (.A(sr_new[8]), .B(\inf_abs1_a_2[8] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[8] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I3_P0N (.A(sum_3), .B(
        \un1_next_sum[0] ), .Y(N481));
    AO1 next_ireg_3_0_ADD_22x22_fast_I76_Y (.A(N349), .B(N346), .C(
        N345), .Y(N384));
    DFN1E1C0 \sumreg[21]  (.D(\next_sum[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_21));
    NOR3B \ireg_RNI2M741[11]  (.A(\state[3]_net_1 ), .B(
        \ireg[11]_net_1 ), .C(integral_1_0), .Y(\ireg_m[11] ));
    OR3 \ireg_RNI869D2[25]  (.A(\un3_next_sum_m[25] ), .B(
        \un1_next_sum_0_iv_0[25] ), .C(\ireg_m[25] ), .Y(
        \un1_next_sum_0_iv[25] ));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I143_un1_Y (.A(N407), .B(N423), 
        .C(N359), .Y(I143_un1_Y));
    MX2 \p_adj_RNO[7]  (.A(sr_new[7]), .B(\inf_abs1_a_2[7] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[7] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I84_Y (.A(N516), .B(N520), .C(
        N519), .Y(N634));
    AO1 next_ireg_3_0_ADD_22x22_fast_I42_Y (.A(N284), .B(N288), .C(
        N287), .Y(N347));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I222_Y (.A(I222_un1_Y), .B(N699), 
        .Y(N781));
    XA1B \sumreg_RNO[36]  (.A(N1027), .B(ADD_40x40_fast_I454_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[36] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I1_P0N (.A(sum_1_d0), .B(
        \un1_next_sum[0] ), .Y(N475));
    OA1 next_ireg_3_0_ADD_22x22_fast_I31_Y (.A(\i_adj[12]_net_1 ), .B(
        \i_adj[14]_net_1 ), .C(N306), .Y(N336));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I380_un1_Y_0 (.A(N874), .B(
        N821), .Y(ADD_40x40_fast_I380_un1_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I129_Y (.A(
        ADD_22x22_fast_I129_un1_Y_0), .B(N531), .C(
        ADD_22x22_fast_I129_Y_0), .Y(N507));
    OR3 next_ireg_3_0_ADD_22x22_fast_I143_Y (.A(I143_un1_Y), .B(
        ADD_22x22_fast_I143_Y_2), .C(I122_un1_Y), .Y(N494));
    DFN1E1C0 \p_adj[1]  (.D(\inf_abs1_5[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[1]_net_1 ));
    NOR3A inf_abs1_a_2_I_27 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .C(
        sr_new[9]), .Y(N_4));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I186_Y (.A(I186_un1_Y), .B(N658), 
        .Y(N739));
    NOR2 inf_abs2_a_0_I_15 (.A(integral[9]), .B(integral[10]), .Y(
        \DWACT_FINC_E[1] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I434_Y_0 (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(ADD_40x40_fast_I434_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I227_Y (.A(N704), .B(N712), .Y(
        N786));
    DFN1E1C0 \p_adj[7]  (.D(\inf_abs1_5[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[7]_net_1 ));
    OR2 \ireg_RNIINPP1[8]  (.A(\un3_next_sum_m[8] ), .B(
        \un1_next_sum_iv_0[8] ), .Y(\un1_next_sum_iv_2[8] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I299_Y (.A(N802), .B(N786), .Y(
        N870));
    DFN1E1C0 \sumreg[11]  (.D(\next_sum[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_11));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I433_Y_0 (.A(sum_15), .B(
        \un1_next_sum[15] ), .Y(ADD_40x40_fast_I433_Y_0));
    NOR3B \preg_RNI7QBI[13]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[13]_net_1 ), .Y(\un24_next_sum_m[13] ));
    XA1B \sumreg_RNO[33]  (.A(N1033), .B(ADD_40x40_fast_I451_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[33] ));
    DFN1E1C0 \ireg[19]  (.D(\next_ireg_3[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[19]_net_1 ));
    MX2 \i_adj_RNO[10]  (.A(integral[16]), .B(\inf_abs2_a_0[10] ), .S(
        integral_1_0), .Y(\inf_abs2_5[10] ));
    XNOR2 inf_abs2_a_0_I_40 (.A(integral[20]), .B(N_13), .Y(
        \inf_abs2_a_0[14] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I385_Y_0 (.A(N693), .B(N686), .C(
        N685), .Y(ADD_40x40_fast_I385_Y_0));
    NOR2B \preg_RNIBUBI_0[17]  (.A(\preg[17]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[17] ));
    AND3 inf_abs2_a_0_I_54 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E[9] ), .C(\DWACT_FINC_E[12] ), .Y(
        \DWACT_FINC_E[13] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I180_Y (.A(N656), .B(N653), .C(
        N652), .Y(N733));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I167_Y (.A(\i_adj[7]_net_1 ), .B(
        \i_adj[9]_net_1 ), .C(N525), .Y(\next_ireg_3[13] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I57_Y (.A(\sumreg[30]_net_1 ), 
        .B(\sumreg[29]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N607)
        );
    DFN1C0 \state[1]  (.D(\state_RNIEBE9[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[1]_net_1 ));
    OR2 \ireg_RNIIJGV1[10]  (.A(\un3_next_sum_m[10] ), .B(
        \un1_next_sum_iv_0[10] ), .Y(\un1_next_sum_iv_2[10] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I382_Y (.A(
        ADD_40x40_fast_I382_Y_1), .B(I382_un1_Y), .C(I338_un1_Y), .Y(
        N1029));
    MX2 \p_adj_RNO[10]  (.A(sr_new[10]), .B(\inf_abs1_a_2[10] ), .S(
        sr_new_1_0), .Y(\inf_abs1_5[10] ));
    DFN1E1C0 \ireg[22]  (.D(\next_ireg_3[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[22]_net_1 ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I20_P0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[20] ), .C(sum_20), .Y(N532));
    AX1D next_ireg_3_0_ADD_22x22_fast_I169_Y (.A(N424), .B(I133_un1_Y), 
        .C(ADD_22x22_fast_I169_Y_0), .Y(\next_ireg_3[15] ));
    NOR3B \ireg_RNI79NI[9]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[9]_net_1 ), .C(integral_0_0), .Y(\ireg_m[9] ));
    NOR3B inf_abs2_a_0_I_16 (.A(\DWACT_FINC_E[1] ), .B(
        \DWACT_FINC_E_0[0] ), .C(integral[11]), .Y(N_21));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I278_un1_Y (.A(N692), .B(N684), 
        .C(N781), .Y(I278_un1_Y));
    NOR3B inf_abs2_a_0_I_55 (.A(\DWACT_FINC_E[13] ), .B(
        \DWACT_FINC_E[28] ), .C(integral[24]), .Y(N_8));
    DFN1E1C0 \preg[13]  (.D(\p_adj[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[13]_net_1 ));
    DFN1E1C0 \i_adj[6]  (.D(\inf_abs2_5[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[6]_net_1 ));
    DFN1E1C0 \i_adj[4]  (.D(\inf_abs2_5[4] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[4]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I63_Y (.A(N332), .B(N336), .Y(
        N371));
    NOR3C un1_sumreg_0_0_ADD_m8_i_a4_0 (.A(ADD_m8_i_a4_0_0), .B(
        sum_2_d0), .C(N_232), .Y(ADD_m8_i_a4_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I230_Y (.A(N715), .B(N708), .C(
        N707), .Y(N789));
    OR2 \ireg_RNIIDVL1[19]  (.A(\un1_next_sum_iv_0[19] ), .B(
        \un1_next_sum_2[4] ), .Y(\un1_next_sum[19] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I81_Y (.A(sum_17), .B(
        \un1_next_sum[17] ), .C(N526), .Y(N631));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I379_Y_2 (.A(N596), .B(
        ADD_40x40_fast_I379_Y_0), .C(N681), .Y(ADD_40x40_fast_I379_Y_2)
        );
    MX2 \i_adj_RNO[18]  (.A(integral[24]), .B(\inf_abs2_a_0[18] ), .S(
        integral_1_0), .Y(\inf_abs2_5[18] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I250_Y (.A(N735), .B(N728), .C(
        N727), .Y(N809));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I142_un1_Y (.A(N618), .B(N615), 
        .Y(I142_un1_Y));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I456_Y_0 (.A(
        \sumreg[38]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I456_Y_0));
    NOR2A inf_abs1_a_2_I_11 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .Y(
        N_10));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I348_Y (.A(I286_un1_Y), .B(N773), 
        .C(I348_un1_Y), .Y(N1043));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I165_Y (.A(N641), .B(N637), .Y(
        N718));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I381_Y_1 (.A(N600), .B(N596), .C(
        N685), .Y(ADD_40x40_fast_I381_Y_1));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I92_Y (.A(N504_0), .B(sum_12), 
        .C(\un1_next_sum[12] ), .Y(N642));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I348_un1_Y (.A(N774), .B(N790), 
        .C(N1091), .Y(I348_un1_Y));
    DFN1E1C0 \i_adj[9]  (.D(\inf_abs2_5[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[9]_net_1 ));
    NOR2A un1_sumreg_0_0_ADD_40x40_fast_I26_G0N (.A(\sumreg[26]_net_1 )
        , .B(\un1_next_sum_1_iv[26] ), .Y(N549));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I85_Y (.A(sum_15), .B(
        \un1_next_sum[15] ), .C(N520), .Y(N635));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I11_G0N (.A(\un1_next_sum[11] )
        , .B(sum_11), .Y(N504_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I201_Y (.A(
        ADD_40x40_fast_I201_Y_0), .B(N686), .Y(N760));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I72_Y (.A(N534), .B(N538), .C(
        N537), .Y(N622));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I0_S (.A(\i_adj[0]_net_1 ), .B(
        \i_adj[2]_net_1 ), .Y(\next_ireg_3[6] ));
    DFN1E1C0 \i_adj[3]  (.D(\inf_abs2_5[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[3]_net_1 ));
    XA1B \sumreg_RNO[15]  (.A(N1085), .B(ADD_40x40_fast_I433_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[15] ));
    OR2 \preg_RNI5E361[12]  (.A(next_sum_0_sqmuxa_1), .B(
        \un24_next_sum_m[12] ), .Y(\un1_next_sum_iv_0[12] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I242_Y (.A(N727), .B(N720), .C(
        N719), .Y(N801));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y_1 (.A(N371), .B(N378), .C(
        ADD_22x22_fast_I126_Y_0), .Y(ADD_22x22_fast_I126_Y_1));
    OA1 next_ireg_3_0_ADD_22x22_fast_I51_Y (.A(\i_adj[3]_net_1 ), .B(
        \i_adj[5]_net_1 ), .C(N273), .Y(N356));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I178_Y (.A(\i_adj[18]_net_1 ), 
        .B(\i_adj[20]_net_1 ), .C(N494), .Y(\next_ireg_3[24] ));
    XA1 \ireg_RNIOGDP[19]  (.A(integral_0_0), .B(\ireg[19]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[19] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I231_Y (.A(N716), .B(N708), .Y(
        N790));
    OR3 \preg_RNIJD562[18]  (.A(\un24_next_sum_m[18] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[18] ), .Y(
        \un1_next_sum_iv_2[18] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I184_Y (.A(N660), .B(N657), .C(
        N656), .Y(N737));
    XNOR2 inf_abs2_a_0_I_56 (.A(integral[25]), .B(N_8), .Y(
        \inf_abs2_a_0[19] ));
    OR3 \preg_RNIKPPP1[9]  (.A(\un24_next_sum_m[9] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[9] ), .Y(
        \un1_next_sum_iv_2[9] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I87_Y (.A(I87_un1_Y), .B(N357), 
        .Y(N396));
    DFN1E1C0 \sumreg[34]  (.D(\next_sum[34] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[34]_net_1 ));
    OR2 \preg_RNI3C4M3[13]  (.A(\un1_next_sum_iv_2[13] ), .B(
        \un1_next_sum_iv_1[13] ), .Y(\un1_next_sum[13] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I340_un1_Y (.A(N848), .B(N879), 
        .Y(I340_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I247_Y (.A(N724), .B(N732), .Y(
        N806));
    DFN1C0 \state_0[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_0[2]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I60_Y (.A(\sumreg[27]_net_1 ), 
        .B(\sumreg[28]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N610)
        );
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I385_un1_Y (.A(N884), .B(
        \un1_next_sum[0] ), .C(N852), .Y(I385_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I173_Y (.A(N645), .B(N649), .Y(
        N726));
    DFN1E1C0 \ireg[7]  (.D(\next_ireg_3[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[7]_net_1 ));
    XA1B \sumreg_RNO[28]  (.A(N1046), .B(ADD_40x40_fast_I446_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[28] ));
    OR2 \state_RNIQM1C1[4]  (.A(N_232), .B(\un1_next_sum_2[4] ), .Y(
        N_228));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I380_un1_Y (.A(N774), .B(N758), 
        .C(ADD_40x40_fast_I380_un1_Y_0), .Y(I380_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I238_Y (.A(N723), .B(N716), .C(
        N715), .Y(N797));
    XA1B \sumreg_RNO[3]  (.A(\un1_next_sum[0] ), .B(
        ADD_40x40_fast_I421_Y_0), .C(\state[2]_net_1 ), .Y(
        \next_sum[3] ));
    DFN1E1C0 \preg[7]  (.D(\p_adj[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[7]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I44_Y (.A(\sumreg[35]_net_1 ), 
        .B(\sumreg[36]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N594)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I258_Y (.A(N736), .B(N743), .C(
        N735), .Y(N817));
    OR3 next_ireg_3_0_ADD_22x22_fast_I131_Y (.A(I131_un1_Y), .B(
        ADD_22x22_fast_I131_Y_0), .C(I106_un1_Y), .Y(N513));
    DFN1E1C0 \ireg[16]  (.D(\next_ireg_3[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[16]_net_1 ));
    NOR2B \state_RNIR7Q8[5]  (.A(\state[5]_net_1 ), .B(sr_new[12]), .Y(
        next_sum_0_sqmuxa_2));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I273_Y (.A(N760), .B(N776), .Y(
        N844));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I195_Y_0 (.A(\sumreg[37]_net_1 )
        , .B(\sumreg[38]_net_1 ), .C(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I195_Y_0));
    XA1B \sumreg_RNO[32]  (.A(N1035), .B(ADD_40x40_fast_I450_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[32] ));
    DFN1E1C0 \preg[10]  (.D(\p_adj[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[10]_net_1 ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I163_Y_0 (.A(\i_adj[3]_net_1 ), 
        .B(\i_adj[5]_net_1 ), .Y(ADD_22x22_fast_I163_Y_0));
    DFN1E1C0 \preg[18]  (.D(\p_adj[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[18]_net_1 ));
    NOR3 inf_abs2_a_0_I_18 (.A(integral[10]), .B(integral[9]), .C(
        integral[11]), .Y(\DWACT_FINC_E[2] ));
    XA1B \sumreg_RNO[8]  (.A(N1106), .B(ADD_40x40_fast_I426_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[8] ));
    NOR3B \ireg_RNI5M101[15]  (.A(integral_0_0), .B(\state[3]_net_1 ), 
        .C(\ireg[15]_net_1 ), .Y(\un3_next_sum_m[15] ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I23_Y (.A(\i_adj[16]_net_1 ), .B(
        \i_adj[18]_net_1 ), .C(N_9), .Y(N328));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I178_Y (.A(N654), .B(N651), .C(
        N650), .Y(N731));
    NOR2B inf_abs2_a_0_I_34 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .Y(N_15));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I98_Y (.A(N495), .B(N499), .C(
        N498), .Y(N648));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I7_P0N (.A(
        \un1_next_sum_iv_1[7] ), .B(\un1_next_sum_iv_2[7] ), .C(sum_7), 
        .Y(N493));
    NOR2 inf_abs2_a_0_I_47 (.A(integral[21]), .B(integral[22]), .Y(
        \DWACT_FINC_E[11] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I89_Y (.A(N511), .B(N514), .Y(
        N639));
    NOR2 inf_abs1_a_2_I_21 (.A(sr_new[6]), .B(sr_new[7]), .Y(
        \DWACT_FINC_E_0[3] ));
    AO1 \preg_RNIBIJM1[13]  (.A(\preg[13]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[13] ), .Y(
        \un1_next_sum_iv_1[13] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I5_G0N (.A(\i_adj[7]_net_1 ), 
        .B(\i_adj[5]_net_1 ), .Y(N281));
    AX1D next_ireg_3_0_ADD_22x22_fast_I176_Y (.A(I126_un1_Y), .B(
        ADD_22x22_fast_I126_Y_1), .C(ADD_22x22_fast_I176_Y_0), .Y(
        \next_ireg_3[22] ));
    NOR3 inf_abs2_a_0_I_8 (.A(integral[7]), .B(integral[6]), .C(
        integral[8]), .Y(N_24));
    XA1B \sumreg_RNO[16]  (.A(N1082), .B(ADD_40x40_fast_I434_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[16] ));
    NOR3B inf_abs2_a_0_I_19 (.A(\DWACT_FINC_E[2] ), .B(
        \DWACT_FINC_E_0[0] ), .C(integral[12]), .Y(N_20));
    NOR3B \ireg_RNIF7DP[10]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[10]_net_1 ), .Y(\un3_next_sum_m[10] ));
    NOR2B \state_RNIEBE9[0]  (.A(sum_enable), .B(sum_rdy), .Y(
        \state_RNIEBE9[0]_net_1 ));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I78_Y (.A(N525_0), .B(sum_19), 
        .C(\un1_next_sum[19] ), .Y(N628));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I132_un1_Y (.A(N423), .B(N359), 
        .Y(I132_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I0_CO1 (.A(\i_adj[0]_net_1 ), 
        .B(\i_adj[2]_net_1 ), .Y(N266));
    OR2A un1_sumreg_0_0_ADD_40x40_fast_I26_P0N (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[26]_net_1 ), .Y(N550));
    OR2 \ireg_RNIHB562[17]  (.A(\un3_next_sum_m[17] ), .B(
        \un1_next_sum_iv_0[17] ), .Y(\un1_next_sum_iv_2[17] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I229_Y (.A(N706), .B(N714), .Y(
        N788));
    XA1B \sumreg_RNO[13]  (.A(N1091), .B(ADD_40x40_fast_I431_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[13] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I112_un1_Y (.A(N387), .B(N394), 
        .Y(I112_un1_Y));
    XNOR2 inf_abs2_a_0_I_7 (.A(integral[8]), .B(N_25), .Y(
        \inf_abs2_a_0[2] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I133_un1_Y (.A(N425), .B(N266), 
        .Y(I133_un1_Y));
    XNOR2 inf_abs2_a_0_I_35 (.A(integral[18]), .B(N_15), .Y(
        \inf_abs2_a_0[12] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I1_P0N (.A(\i_adj[1]_net_1 ), .B(
        \i_adj[3]_net_1 ), .Y(N270));
    XOR2 inf_abs2_a_0_I_5 (.A(integral[6]), .B(integral[7]), .Y(
        \inf_abs2_a_0[1] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I332_un1_Y (.A(N772), .B(N756), 
        .C(N871), .Y(I332_un1_Y));
    AND3 inf_abs2_a_0_I_61 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[15] ), .Y(N_6));
    AND3 inf_abs2_a_0_I_58 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[14] ), .Y(N_7_0));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I111_Y (.A(\un1_next_sum[0] ), 
        .B(sum_2_d0), .C(N481), .Y(N661));
    XA1B \sumreg_RNO[19]  (.A(N1073), .B(ADD_40x40_fast_I437_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[19] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I68_Y (.A(N341), .B(N338), .C(
        N337), .Y(N376));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I16_G0N (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(N519));
    XNOR2 inf_abs1_a_2_I_12 (.A(sr_new[4]), .B(N_10), .Y(
        \inf_abs1_a_2[4] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I446_Y_0 (.A(
        \sumreg[28]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I446_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I109_Y (.A(N391), .B(N383), .Y(
        N423));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I93_Y (.A(sum_12), .B(
        \un1_next_sum[12] ), .C(N505), .Y(N643));
    DFN1E1C0 \p_adj[12]  (.D(\inf_abs1_5[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[12]_net_1 ));
    DFN1E1C0 \p_adj[2]  (.D(\inf_abs1_5[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[2]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I138_un1_Y (.A(N614), .B(N611), 
        .Y(I138_un1_Y));
    MX2 \i_adj_RNO[9]  (.A(integral[15]), .B(\inf_abs2_a_0[9] ), .S(
        integral[25]), .Y(\inf_abs2_5[9] ));
    DFN1E1C0 \ireg[18]  (.D(\next_ireg_3[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[18]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_1 (.A(N328), .B(N331), .C(
        ADD_22x22_fast_I143_Y_0), .Y(ADD_22x22_fast_I143_Y_1));
    NOR3A inf_abs2_a_0_I_13 (.A(\DWACT_FINC_E_0[0] ), .B(integral[9]), 
        .C(integral[10]), .Y(N_22));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I313_Y (.A(N816), .B(N800), .Y(
        N884));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I73_Y (.A(sum_21), .B(
        \un1_next_sum[21] ), .C(N538), .Y(N623));
    NOR3B \ireg_RNI68NI[8]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[8]_net_1 ), .C(integral_0_0), .Y(\ireg_m[8] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I45_Y (.A(\sumreg[36]_net_1 ), 
        .B(\sumreg[35]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N595)
        );
    NOR2B \preg_RNIATBI_0[16]  (.A(\preg[16]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[16] ));
    DFN1E1C0 \ireg[9]  (.D(\next_ireg_3[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[9]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I382_Y_0 (.A(N679), .B(N687), .Y(
        ADD_40x40_fast_I382_Y_0));
    DFN1E1C0 \preg[14]  (.D(\p_adj[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[14]_net_1 ));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I96_Y (.A(N498), .B(sum_10), .C(
        \un1_next_sum[10] ), .Y(N646));
    XNOR2 inf_abs2_a_0_I_59 (.A(integral[25]), .B(N_7_0), .Y(
        \inf_abs2_a_0[20] ));
    AND3 inf_abs2_a_0_I_24 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E_0[4] ));
    DFN1E1C0 \preg[9]  (.D(\p_adj[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[9]_net_1 ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I426_Y_0 (.A(sum_8), .B(
        \un1_next_sum[8] ), .Y(ADD_40x40_fast_I426_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I379_Y (.A(
        ADD_40x40_fast_I379_un1_Y_0), .B(N819), .C(
        ADD_40x40_fast_I379_Y_4), .Y(N1023));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I222_un1_Y (.A(N707), .B(N700), 
        .Y(I222_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I76_Y (.A(N528_0), .B(N532), .C(
        N531_0), .Y(N626));
    DFN1P0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .PRE(n_rst_c), 
        .Q(sum_rdy));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I205_Y (.A(N682), .B(N690), .Y(
        N764));
    NOR2B inf_abs1_a_2_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_2));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I177_Y (.A(N649), .B(N653), .Y(
        N730));
    NOR3B inf_abs2_a_0_I_36 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .C(integral[18]), .Y(N_14));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I8_G0N (.A(\un1_next_sum[8] ), 
        .B(sum_8), .Y(N495));
    XA1B \sumreg_RNO[6]  (.A(N819), .B(ADD_40x40_fast_I424_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[6] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I218_un1_Y (.A(N619), .B(N615), 
        .C(N703), .Y(I218_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I71_Y (.A(N344), .B(N340), .Y(
        N379));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I145_Y (.A(N621), .B(N617), .Y(
        N698));
    AO1A \state_RNO[0]  (.A(sum_enable), .B(sum_rdy), .C(
        \state[5]_net_1 ), .Y(\state_ns[0] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I62_Y (.A(\sumreg[26]_net_1 ), 
        .B(\sumreg[27]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N612)
        );
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I380_Y (.A(I380_un1_Y), .B(
        ADD_40x40_fast_I380_Y_2), .C(I334_un1_Y), .Y(N1025));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I235_Y (.A(N720), .B(N712), .Y(
        N794));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I191_Y (.A(N664), .B(I116_un1_Y), 
        .Y(N745));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I455_Y_0 (.A(
        \sumreg[37]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I455_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I255_Y (.A(N740), .B(N732), .Y(
        N814));
    AO1 next_ireg_3_0_ADD_22x22_fast_I82_Y (.A(N355), .B(N352), .C(
        N351), .Y(N390));
    NOR2A inf_abs2_a_0_I_25 (.A(\DWACT_FINC_E_0[4] ), .B(integral[14]), 
        .Y(N_18));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I183_Y (.A(N484), .B(N481), .C(
        N655), .Y(N736));
    DFN1E1C0 \ireg[8]  (.D(\next_ireg_3[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[8]_net_1 ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I25_Y (.A(\i_adj[16]_net_1 ), .B(
        \i_adj[18]_net_1 ), .C(N312), .Y(N330));
    OA1 next_ireg_3_0_ADD_22x22_fast_I43_Y (.A(\i_adj[6]_net_1 ), .B(
        \i_adj[8]_net_1 ), .C(N288), .Y(N348));
    XNOR2 inf_abs1_a_2_I_35 (.A(sr_new[12]), .B(N_2), .Y(
        \inf_abs1_a_2[12] ));
    DFN1E1C0 \preg[8]  (.D(\p_adj[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[8]_net_1 ));
    XNOR2 inf_abs2_a_0_I_53 (.A(integral[24]), .B(N_9_0), .Y(
        \inf_abs2_a_0[18] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I301_Y (.A(N804), .B(N788), .Y(
        N872));
    DFN1E1C0 \i_adj[14]  (.D(\inf_abs2_5[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[14]_net_1 ));
    NOR3B \preg_RNIBKDK[8]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[8]_net_1 ), .Y(\un24_next_sum_m[8] ));
    DFN1E1C0 \sumreg[32]  (.D(\next_sum[32] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[32]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I108_un1_Y (.A(N480), .B(N484), 
        .Y(I108_un1_Y));
    AO1 \preg_RNI1P241[8]  (.A(\preg[8]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[8] ), .Y(
        \un1_next_sum_iv_1[8] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I346_Y (.A(
        ADD_40x40_fast_I346_un1_Y_0), .B(N1085), .C(
        ADD_40x40_fast_I346_Y_0), .Y(N1037));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I28_Y (.A(N305), .B(
        \i_adj[16]_net_1 ), .C(\i_adj[14]_net_1 ), .Y(N333));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I249_Y (.A(N726), .B(N734), .Y(
        N808));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I351_Y (.A(I292_un1_Y), .B(N779), 
        .C(I351_un1_Y), .Y(N1052));
    MX2 \i_adj_RNO[6]  (.A(integral[12]), .B(\inf_abs2_a_0[6] ), .S(
        integral_1_0), .Y(\inf_abs2_5[6] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I188_Y (.A(N664), .B(N661), .C(
        N660), .Y(N741));
    AND3 inf_abs1_a_2_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(N_6_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I16_P0N (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(N520));
    NOR3B \preg_RNICVBI[18]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[18]_net_1 ), .Y(\un24_next_sum_m[18] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I49_Y (.A(\sumreg[34]_net_1 ), 
        .B(\sumreg[33]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N599)
        );
    XNOR2 inf_abs2_a_0_I_26 (.A(integral[15]), .B(N_18), .Y(
        \inf_abs2_a_0[9] ));
    XA1B \sumreg_RNO[12]  (.A(N1094), .B(ADD_40x40_fast_I430_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[12] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I54_Y (.A(\sumreg[31]_net_1 ), 
        .B(\sumreg[30]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N604)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I315_Y (.A(N804), .B(N819), .C(
        N803), .Y(N1088));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I112_Y (.A(sum_2_d0), .B(
        sum_1_d0), .C(\un1_next_sum[0] ), .Y(N662));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I177_Y_0 (.A(\i_adj[19]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(ADD_22x22_fast_I177_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I106_Y (.A(N483), .B(N487), .C(
        N486), .Y(N656));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I7_G0N (.A(
        \un1_next_sum_iv_1[7] ), .B(\un1_next_sum_iv_2[7] ), .C(sum_7), 
        .Y(N492_0));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I164_Y (.A(
        ADD_22x22_fast_I164_Y_0), .B(N394), .Y(\next_ireg_3[10] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_1 (.A(
        ADD_22x22_fast_I142_Y_0_a3_0), .B(N329), .C(
        ADD_22x22_fast_I142_Y_0_0), .Y(ADD_22x22_fast_I142_Y_0_1));
    XNOR2 inf_abs2_a_0_I_62 (.A(integral[25]), .B(N_6), .Y(
        \inf_abs2_a_0[21] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I419_Y_0 (.A(sum_1_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I419_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I68_Y (.A(N540), .B(N544), .C(
        N543), .Y(N618));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I22_G0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[22] ), .C(sum_22), .Y(N537));
    NOR2 inf_abs2_a_0_I_38 (.A(integral[18]), .B(integral[19]), .Y(
        \DWACT_FINC_E[8] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I380_Y_2 (.A(N758), .B(N773), .C(
        ADD_40x40_fast_I380_Y_1), .Y(ADD_40x40_fast_I380_Y_2));
    NOR3 inf_abs2_a_0_I_41 (.A(integral[19]), .B(integral[18]), .C(
        integral[20]), .Y(\DWACT_FINC_E[9] ));
    MX2 \p_adj_RNO[9]  (.A(sr_new[9]), .B(\inf_abs1_a_2[9] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[9] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I162_Y_0 (.A(\i_adj[2]_net_1 ), 
        .B(\i_adj[4]_net_1 ), .Y(ADD_22x22_fast_I162_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I136_Y (.A(N612), .B(N608), .Y(
        N689));
    XA1 \ireg_RNI35NI[5]  (.A(integral_0_0), .B(\ireg[5]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[5] ));
    DFN1E1C0 \sumreg[33]  (.D(\next_sum[33] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[33]_net_1 ));
    AO1 \ireg_RNI5LMA1[18]  (.A(\ireg[18]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[18] ), .Y(
        \un1_next_sum_iv_1[18] ));
    XA1B \sumreg_RNO[2]  (.A(N745), .B(ADD_40x40_fast_I420_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[2] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I156_Y (.A(N632), .B(N629), .C(
        N628), .Y(N709));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I352_un1_Y_0 (.A(N798), .B(
        N782), .Y(ADD_40x40_fast_I352_un1_Y_0));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I100_Y (.A(N492_0), .B(sum_8), 
        .C(\un1_next_sum[8] ), .Y(N650));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I165_Y_0 (.A(\i_adj[5]_net_1 ), 
        .B(\i_adj[7]_net_1 ), .Y(ADD_22x22_fast_I165_Y_0));
    DFN1E1C0 \i_adj[12]  (.D(\inf_abs2_5[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[12]_net_1 ));
    NOR3B \ireg_RNI9FKH[9]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[9]_net_1 ), .Y(\un3_next_sum_m[9] ));
    NOR2B \i_adj_RNO[19]  (.A(\inf_abs2_a_0[19] ), .B(integral[25]), 
        .Y(\inf_abs2_5[19] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I39_Y (.A(N291), .B(N294), .Y(
        N344));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y_0 (.A(N335), .B(N332), .C(
        N331), .Y(ADD_22x22_fast_I126_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I14_G0N (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .Y(N308));
    DFN1E1C0 \sumreg[30]  (.D(\next_sum[30] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[30]_net_1 ));
    AND3 inf_abs2_a_0_I_39 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E_0[7] ), .C(\DWACT_FINC_E[8] ), .Y(N_13));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I24_Y (.A(N311), .B(
        \i_adj[16]_net_1 ), .C(\i_adj[18]_net_1 ), .Y(N329));
    OA1 next_ireg_3_0_ADD_22x22_fast_I37_Y (.A(\i_adj[10]_net_1 ), .B(
        \i_adj[12]_net_1 ), .C(N294), .Y(N342));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I302_Y (.A(N805), .B(N790), .C(
        N789), .Y(N873));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I292_un1_Y (.A(N795), .B(N780), 
        .Y(I292_un1_Y));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I130_Y (.A(N606), .B(N602), .Y(
        N683));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I80_Y (.A(N522), .B(N526), .C(
        N525_0), .Y(N630));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I346_un1_Y_0 (.A(N786), .B(
        N770), .Y(ADD_40x40_fast_I346_un1_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I288_un1_Y (.A(N791), .B(N776), 
        .Y(I288_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I0_G0N (.A(N_228), .B(sum_0_d0)
        , .Y(N471));
    NOR3 \state_RNINAIE[6]  (.A(sum_rdy), .B(\state[6]_net_1 ), .C(
        \state_0[1]_net_1 ), .Y(N_416_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I150_Y (.A(N626), .B(N623), .C(
        N622), .Y(N703));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I161_Y (.A(N633), .B(N637), .Y(
        N714));
    AO1 next_ireg_3_0_ADD_22x22_fast_I40_Y (.A(N287), .B(N291), .C(
        N290), .Y(N345));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I346_Y_0 (.A(N785), .B(N770), .C(
        N769), .Y(ADD_40x40_fast_I346_Y_0));
    OA1A un1_sumreg_0_0_ADD_40x40_fast_I63_Y (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[27]_net_1 ), .C(N550), .Y(
        N613));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I187_Y (.A(N484), .B(N481), .C(
        ADD_40x40_fast_I187_Y_0), .Y(N740));
    XA1B \sumreg_RNO[4]  (.A(N823), .B(ADD_40x40_fast_I422_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[4] ));
    OR3 \preg_RNIQRGV1[14]  (.A(\un24_next_sum_m[14] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[14] ), .Y(
        \un1_next_sum_iv_2[14] ));
    NOR2B \state_RNIFFD8[3]  (.A(\state[3]_net_1 ), .B(integral[25]), 
        .Y(next_sum_0_sqmuxa));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I352_Y (.A(
        ADD_40x40_fast_I352_un1_Y_0), .B(N1103), .C(
        ADD_40x40_fast_I352_Y_0), .Y(N1055));
    XA1B \sumreg_RNO[5]  (.A(N821), .B(ADD_40x40_fast_I423_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[5] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I378_Y (.A(
        ADD_40x40_fast_I378_Y_3), .B(I378_un1_Y), .C(I330_un1_Y), .Y(
        N1021));
    OA1 next_ireg_3_0_ADD_22x22_fast_I45_Y (.A(\i_adj[6]_net_1 ), .B(
        \i_adj[8]_net_1 ), .C(N282), .Y(N350));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I171_Y (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .C(N513), .Y(\next_ireg_3[17] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_o3_0_0 (.A(N337), .B(
        N334), .C(N333), .Y(ADD_22x22_fast_I142_Y_0_o3_0_0));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I432_Y_0 (.A(sum_14), .B(
        \un1_next_sum[14] ), .Y(ADD_40x40_fast_I432_Y_0));
    DFN1E1C0 \sumreg[37]  (.D(\next_sum[37] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[37]_net_1 ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I51_Y (.A(\sumreg[33]_net_1 ), 
        .B(\sumreg[32]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N601)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I383_Y_1 (.A(N764), .B(N779), .C(
        ADD_40x40_fast_I383_Y_0), .Y(ADD_40x40_fast_I383_Y_1));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I23_P0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[23] ), .C(sum_23), .Y(N541));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_2 (.A(N367), .B(N374), .C(
        ADD_22x22_fast_I143_Y_1), .Y(ADD_22x22_fast_I143_Y_2));
    AO13 un1_sumreg_0_0_ADD_40x40_fast_I66_Y (.A(\sumreg[25]_net_1 ), 
        .B(N543), .C(\un1_next_sum_0_iv[25] ), .Y(N616));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I445_Y_0 (.A(
        \sumreg[27]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I445_Y_0));
    XNOR2 inf_abs2_a_0_I_28 (.A(integral[16]), .B(N_17), .Y(
        \inf_abs2_a_0[10] ));
    NOR3 inf_abs2_a_0_I_33 (.A(integral[16]), .B(integral[15]), .C(
        integral[17]), .Y(\DWACT_FINC_E_0[7] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I55_Y (.A(\sumreg[30]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N605)
        );
    DFN1C0 \state_1[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_1[2]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I48_Y (.A(N275), .B(N279), .C(
        N278), .Y(N353));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I3_G0N (.A(sum_3), .B(
        \un1_next_sum[0] ), .Y(N480));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I344_un1_Y (.A(N852), .B(N883), 
        .Y(I344_un1_Y));
    MX2 \i_adj_RNO[4]  (.A(integral[10]), .B(\inf_abs2_a_0[4] ), .S(
        integral_1_0), .Y(\inf_abs2_5[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I210_Y (.A(N695), .B(N688), .C(
        N687), .Y(N769));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I15_G0N (.A(\un1_next_sum[15] )
        , .B(sum_15), .Y(N516));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I425_Y_0 (.A(
        \un1_next_sum_iv_1[7] ), .B(\un1_next_sum_iv_2[7] ), .C(sum_7), 
        .Y(ADD_40x40_fast_I425_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I139_Y (.A(N611), .B(N615), .Y(
        N692));
    OR2B next_ireg_3_0_ADD_22x22_fast_I17_G0N_i (.A(\i_adj[19]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(N_7));
    XA1 \ireg_RNIKDEP[24]  (.A(integral_0_0), .B(\ireg[24]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[24] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I384_un1_Y (.A(N882), .B(N666), 
        .C(N850), .Y(I384_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I277_Y (.A(N764), .B(N780), .Y(
        N848));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I159_Y (.A(N635), .B(N631), .Y(
        N712));
    DFN1E1C0 \i_adj[13]  (.D(\inf_abs2_5[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[13]_net_1 ));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I104_Y (.A(N486), .B(sum_6), .C(
        \un1_next_sum[6] ), .Y(N654));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I115_un1_Y (.A(N393), .B(N266), 
        .Y(I115_un1_Y));
    NOR3 inf_abs2_a_0_I_29 (.A(integral[14]), .B(integral[13]), .C(
        integral[12]), .Y(\DWACT_FINC_E[5] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I130_Y_0 (.A(N386), .B(N379), .C(
        N378), .Y(ADD_22x22_fast_I130_Y_0));
    DFN1E1C0 \preg[12]  (.D(\p_adj[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[12]_net_1 ));
    MX2 \i_adj_RNO[2]  (.A(integral[8]), .B(\inf_abs2_a_0[2] ), .S(
        integral_1_0), .Y(\inf_abs2_5[2] ));
    DFN1E1C0 \i_adj[5]  (.D(\inf_abs2_5[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[5]_net_1 ));
    DFN1E1C0 \ireg[20]  (.D(\next_ireg_3[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[20]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I379_Y_0 (.A(\sumreg[36]_net_1 )
        , .B(\sumreg[37]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(
        ADD_40x40_fast_I379_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I321_un1_Y (.A(N816), .B(
        \un1_next_sum[0] ), .Y(I321_un1_Y));
    OR3 un1_sumreg_0_0_ADD_m8_i_o4_1 (.A(sum_2_d0), .B(sum_1_d0), .C(
        sum_0_d0), .Y(ADD_m8_i_o4_1));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I378_Y_0 (.A(\sumreg[38]_net_1 )
        , .B(\sumreg[37]_net_1 ), .C(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I378_Y_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I2_P0N (.A(\i_adj[2]_net_1 ), .B(
        \i_adj[4]_net_1 ), .Y(N273));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I134_Y (.A(N610), .B(N606), .Y(
        N687));
    DFN1E1C0 \i_adj[0]  (.D(\inf_abs2_5[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[0]_net_1 ));
    DFN1E1C0 \p_adj[6]  (.D(\inf_abs1_5[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[6]_net_1 ));
    MX2 \p_adj_RNO[4]  (.A(sr_new[4]), .B(\inf_abs1_a_2[4] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I154_Y (.A(N630), .B(N627), .C(
        N626), .Y(N707));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I211_Y (.A(N619), .B(N615), .C(
        N688), .Y(N770));
    AO1A \ireg_RNIOTDU1[12]  (.A(\ireg[12]_net_1 ), .B(
        next_sum_0_sqmuxa), .C(\un1_next_sum_iv_0[12] ), .Y(
        \un1_next_sum_iv_2[12] ));
    NOR3B \ireg_RNI46NI[6]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[6]_net_1 ), .C(integral_0_0), .Y(\ireg_m[6] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I12_G0N (.A(\un1_next_sum[12] )
        , .B(sum_12), .Y(N507_0));
    XA1B \sumreg_RNO[24]  (.A(N1058), .B(ADD_40x40_fast_I442_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[24] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I59_Y (.A(N328), .B(N332), .Y(
        N367));
    MX2 \i_adj_RNO[0]  (.A(integral[6]), .B(integral[6]), .S(
        integral_1_0), .Y(\inf_abs2_5[0] ));
    AND3 inf_abs2_a_0_I_42 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E_0[7] ), .C(\DWACT_FINC_E[9] ), .Y(N_12_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I17_P0N_i_o3 (.A(
        \i_adj[19]_net_1 ), .B(\i_adj[17]_net_1 ), .Y(N_9));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I218_Y (.A(I218_un1_Y), .B(N695), 
        .Y(N777));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I168_Y_0 (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[8]_net_1 ), .Y(ADD_22x22_fast_I168_Y_0));
    XNOR2 inf_abs2_a_0_I_23 (.A(integral[14]), .B(N_19), .Y(
        \inf_abs2_a_0[8] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I66_Y (.A(N339), .B(N336), .C(
        N335), .Y(N374));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I44_Y (.A(N281), .B(
        \i_adj[6]_net_1 ), .C(\i_adj[8]_net_1 ), .Y(N349));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I439_Y_0 (.A(sum_21), .B(
        \un1_next_sum[21] ), .Y(ADD_40x40_fast_I439_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I450_Y_0 (.A(
        \sumreg[32]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I450_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I234_Y (.A(N719), .B(N712), .C(
        N711), .Y(N793));
    NOR3 inf_abs1_a_2_I_33 (.A(sr_new[10]), .B(sr_new[9]), .C(
        sr_new[11]), .Y(\DWACT_FINC_E[7] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I384_Y (.A(N850), .B(N881), .C(
        ADD_40x40_fast_I384_Y_2), .Y(N1033));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I254_Y (.A(N739), .B(N732), .C(
        N731), .Y(N813));
    MX2 \i_adj_RNO[7]  (.A(integral[13]), .B(\inf_abs2_a_0[7] ), .S(
        integral[25]), .Y(\inf_abs2_5[7] ));
    DFN1E1C0 \i_adj[21]  (.D(\inf_abs2_5[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[21]_net_1 ));
    XA1B \sumreg_RNO[9]  (.A(N1103), .B(ADD_40x40_fast_I427_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[9] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I59_Y (.A(\sumreg[28]_net_1 ), 
        .B(\sumreg[29]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N609)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I162_Y (.A(N638), .B(N635), .C(
        N634), .Y(N715));
    NOR3B \ireg_RNI7DKH[7]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[7]_net_1 ), .Y(\un3_next_sum_m[7] ));
    AO1 \ireg_RNI3JMA1[17]  (.A(\ireg[17]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[17] ), .Y(
        \un1_next_sum_iv_1[17] ));
    DFN1E1C0 \ireg[14]  (.D(\next_ireg_3[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[14]_net_1 ));
    OR2 \preg_RNIR34M3[11]  (.A(\un1_next_sum_iv_2[11] ), .B(
        \un1_next_sum_iv_1[11] ), .Y(\un1_next_sum[11] ));
    DFN1E1C0 \p_adj[11]  (.D(\inf_abs1_5[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[11]_net_1 ));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I82_Y (.A(N519), .B(sum_17), .C(
        \un1_next_sum[17] ), .Y(N632));
    DFN1E1C0 \i_adj[16]  (.D(\inf_abs2_5[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[16]_net_1 ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I4_P0N (.A(\i_adj[6]_net_1 ), .B(
        \i_adj[4]_net_1 ), .Y(N279));
    AO1 next_ireg_3_0_ADD_22x22_fast_I131_Y_0 (.A(N345), .B(N342), .C(
        N341), .Y(ADD_22x22_fast_I131_Y_0));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I437_Y_0 (.A(sum_19), .B(
        \un1_next_sum[19] ), .Y(ADD_40x40_fast_I437_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I268_un1_Y (.A(N756), .B(N771), 
        .Y(I268_un1_Y));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I13_P0N (.A(\un1_next_sum[13] ), 
        .B(sum_13), .Y(N511));
    AO1 \ireg_RNIVEMA1[15]  (.A(\ireg[15]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[15] ), .Y(
        \un1_next_sum_iv_1[15] ));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I32_Y (.A(N299), .B(
        \i_adj[12]_net_1 ), .C(\i_adj[14]_net_1 ), .Y(N337));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I352_Y_0 (.A(N797), .B(N782), .C(
        N781), .Y(ADD_40x40_fast_I352_Y_0));
    MX2 \i_adj_RNO[11]  (.A(integral[17]), .B(\inf_abs2_a_0[11] ), .S(
        integral_1_0), .Y(\inf_abs2_5[11] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I130_un1_Y_0 (.A(N387), .B(N379)
        , .Y(ADD_22x22_fast_I130_un1_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I15_G0N (.A(\i_adj[17]_net_1 ), 
        .B(\i_adj[15]_net_1 ), .Y(N311));
    NOR3B \ireg_RNI1L741[10]  (.A(\state[3]_net_1 ), .B(
        \ireg[10]_net_1 ), .C(integral_1_0), .Y(\ireg_m[10] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I298_Y (.A(N801), .B(N786), .C(
        N785), .Y(N869));
    DFN1E1C0 \ireg[4]  (.D(\i_adj[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[4]_net_1 ));
    MX2 \p_adj_RNO[11]  (.A(sr_new[11]), .B(\inf_abs1_a_2[11] ), .S(
        sr_new_1_0), .Y(\inf_abs1_5[11] ));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I172_Y (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[12]_net_1 ), .C(N510), .Y(\next_ireg_3[18] ));
    XA1B \sumreg_RNO[37]  (.A(N1025), .B(ADD_40x40_fast_I455_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[37] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I381_un1_Y (.A(N876), .B(N823), 
        .C(N844), .Y(I381_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I141_Y (.A(N613), .B(N617), .Y(
        N694));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I83_Y (.A(N356), .B(N352), .Y(
        N391));
    AO1 \preg_RNI5CJM1[10]  (.A(\preg[10]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[10] ), .Y(
        \un1_next_sum_iv_1[10] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I111_Y (.A(N393), .B(N385), .Y(
        N425));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I175_Y (.A(N647), .B(N651), .Y(
        N728));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I378_un1_Y_0 (.A(N870), .B(
        N817), .Y(ADD_40x40_fast_I378_un1_Y_0));
    NOR3B \ireg_RNI4O741[13]  (.A(\state[3]_net_1 ), .B(
        \ireg[13]_net_1 ), .C(integral_1_0), .Y(\ireg_m[13] ));
    DFN1E1C0 \sumreg[24]  (.D(\next_sum[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(\sumreg[24]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I26_Y (.A(N308), .B(N312), .C(
        N311), .Y(N331));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I24_G0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[24] ), .C(\sumreg[24]_net_1 ), .Y(N543));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I175_Y (.A(\i_adj[17]_net_1 ), 
        .B(\i_adj[15]_net_1 ), .C(N_11), .Y(\next_ireg_3[21] ));
    NOR3B \ireg_RNI7O101[17]  (.A(integral_0_0), .B(\state[3]_net_1 ), 
        .C(\ireg[17]_net_1 ), .Y(\un3_next_sum_m[17] ));
    AO1 \ireg_RNITCMA1[14]  (.A(\ireg[14]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[14] ), .Y(
        \un1_next_sum_iv_1[14] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I431_Y_0 (.A(sum_13), .B(
        \un1_next_sum[13] ), .Y(ADD_40x40_fast_I431_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I300_Y (.A(N803), .B(N788), .C(
        N787), .Y(N871));
    NOR3B \preg_RNI9SBI[15]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[15]_net_1 ), .Y(\un24_next_sum_m[15] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I103_Y (.A(sum_6), .B(
        \un1_next_sum[6] ), .C(N493), .Y(N653));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I88_Y (.A(N510_0), .B(N514), .C(
        N513_0), .Y(N638));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I0_P0N (.A(N_228), .B(sum_0_d0), 
        .Y(N472));
    NOR3B un1_sumreg_0_0_ADD_40x40_fast_I64_un1_Y (.A(
        \sumreg[25]_net_1 ), .B(N550), .C(\un1_next_sum_0_iv[25] ), .Y(
        I64_un1_Y));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I260_Y (.A(I260_un1_Y), .B(N739), 
        .Y(N821));
    NOR2B \preg_RNI9SBI_0[15]  (.A(\preg[15]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[15] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I379_un1_Y_0 (.A(N772), .B(
        N756), .C(N872), .Y(ADD_40x40_fast_I379_un1_Y_0));
    MX2 \i_adj_RNO[15]  (.A(integral[21]), .B(\inf_abs2_a_0[15] ), .S(
        integral_1_0), .Y(\inf_abs2_5[15] ));
    DFN1E1C0 \sumreg[14]  (.D(\next_sum[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_14));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I350_Y (.A(I290_un1_Y), .B(N777), 
        .C(I350_un1_Y), .Y(N1049));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I203_Y (.A(N680), .B(N688), .Y(
        N762));
    NOR2B \i_adj_RNO[20]  (.A(\inf_abs2_a_0[20] ), .B(integral[25]), 
        .Y(\inf_abs2_5[20] ));
    XNOR2 inf_abs1_a_2_I_14 (.A(sr_new[5]), .B(N_9_1), .Y(
        \inf_abs1_a_2[5] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I170_Y_0 (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[12]_net_1 ), .Y(ADD_22x22_fast_I170_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I133_Y (.A(N605), .B(N609), .Y(
        N686));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I215_Y (.A(N692), .B(N700), .Y(
        N774));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I279_Y (.A(N692), .B(N684), .C(
        N782), .Y(N850));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I153_Y (.A(N625), .B(N629), .Y(
        N706));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I79_Y (.A(N352), .B(N348), .Y(
        N387));
    XA1B \sumreg_RNO[30]  (.A(N1040), .B(ADD_40x40_fast_I448_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[30] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I77_Y (.A(N346), .B(N350), .Y(
        N385));
    XNOR2 inf_abs2_a_0_I_9 (.A(integral[9]), .B(N_24), .Y(
        \inf_abs2_a_0[3] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I233_Y (.A(N718), .B(N710), .Y(
        N792));
    XA1B \sumreg_RNO[31]  (.A(N1037), .B(ADD_40x40_fast_I449_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[31] ));
    NOR3 inf_abs2_a_0_I_10 (.A(integral[7]), .B(integral[6]), .C(
        integral[8]), .Y(\DWACT_FINC_E_0[0] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I440_Y_0 (.A(
        \un1_next_sum_2[4] ), .B(\un1_next_sum_iv_0[22] ), .C(sum_22), 
        .Y(ADD_40x40_fast_I440_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I253_Y (.A(N738), .B(N730), .Y(
        N812));
    AO1 next_ireg_3_0_ADD_22x22_fast_I52_Y (.A(N269), .B(N273), .C(
        N272), .Y(N357));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I108_Y (.A(I108_un1_Y), .B(N483), 
        .Y(N658));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I261_Y (.A(N741), .B(I116_un1_Y), 
        .Y(N823));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I173_Y (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[13]_net_1 ), .C(N507), .Y(\next_ireg_3[19] ));
    NOR3B \preg_RNI9IDK[6]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[6]_net_1 ), .Y(\un24_next_sum_m[6] ));
    NOR2 inf_abs1_a_2_I_15 (.A(sr_new[3]), .B(sr_new[4]), .Y(
        \DWACT_FINC_E_0[1] ));
    XA1B \state_RNIMF7CI9[2]  (.A(N1021), .B(ADD_40x40_fast_I457_Y_0), 
        .C(\state[2]_net_1 ), .Y(\next_sum[39] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I83_Y (.A(sum_17), .B(
        \un1_next_sum[17] ), .C(N520), .Y(N633));
    XA1B \sumreg_RNO[25]  (.A(N1055), .B(ADD_40x40_fast_I443_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[25] ));
    DFN1E1C0 \i_adj[11]  (.D(\inf_abs2_5[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[11]_net_1 ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I307_Y (.A(N728), .B(N736), .C(
        N794), .Y(N878));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I138_Y (.A(I138_un1_Y), .B(N610), 
        .Y(N691));
    DFN1E1C0 \ireg[11]  (.D(\next_ireg_3[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[11]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I311_Y (.A(N814), .B(N798), .Y(
        N882));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I420_Y_0 (.A(sum_2_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I420_Y_0));
    DFN1C0 \state[3]  (.D(\state[6]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[3]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I158_Y (.A(N634), .B(N631), .C(
        N630), .Y(N711));
    MX2 \i_adj_RNO[17]  (.A(integral[23]), .B(\inf_abs2_a_0[17] ), .S(
        integral_1_0), .Y(\inf_abs2_5[17] ));
    DFN1E1C0 \i_adj[1]  (.D(\inf_abs2_5[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[1]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I80_Y (.A(N353), .B(N350), .C(
        N349), .Y(N388));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I86_Y (.A(N513_0), .B(sum_15), 
        .C(\un1_next_sum[15] ), .Y(N636));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I236_Y (.A(N721), .B(N714), .C(
        N713), .Y(N795));
    DFN1E1C0 \sumreg[3]  (.D(\next_sum[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416), .Q(sum_3));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I220_Y (.A(N705), .B(N698), .C(
        N697), .Y(N779));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I256_Y (.A(N741), .B(N734), .C(
        N733), .Y(N815));
    DFN1E1C0 \sumreg_1[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(sum_1_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I382_Y_1 (.A(N762), .B(N777), .C(
        ADD_40x40_fast_I382_Y_0), .Y(ADD_40x40_fast_I382_Y_1));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I4_G0N (.A(\i_adj[6]_net_1 ), 
        .B(\i_adj[4]_net_1 ), .Y(N278));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I357_Y (.A(N876), .B(N823), .C(
        N875), .Y(N1070));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I85_Y (.A(N358), .B(N354), .Y(
        N393));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I24_P0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[24] ), .C(\sumreg[24]_net_1 ), .Y(N544));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I142_Y (.A(I142_un1_Y), .B(N614), 
        .Y(N695));
    DFN1C0 \state_0[1]  (.D(\state_RNIEBE9[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_0[1]_net_1 ));
    NOR3 inf_abs2_a_0_I_50 (.A(integral[22]), .B(integral[21]), .C(
        integral[23]), .Y(\DWACT_FINC_E[12] ));
    NOR3B \preg_RNIAJDK[7]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), .C(
        \preg[7]_net_1 ), .Y(\un24_next_sum_m[7] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I3_G0N (.A(\i_adj[5]_net_1 ), 
        .B(\i_adj[3]_net_1 ), .Y(N275));
    XNOR2 inf_abs1_a_2_I_9 (.A(sr_new[3]), .B(N_11_1), .Y(
        \inf_abs1_a_2[3] ));
    NOR3B inf_abs1_a_2_I_16 (.A(\DWACT_FINC_E_0[1] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[5]), .Y(N_8_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I46_Y (.A(N278), .B(N282), .C(
        N281), .Y(N351));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I13_G0N (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[13]_net_1 ), .Y(N305));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I361_un1_Y (.A(N884), .B(
        \un1_next_sum[0] ), .Y(I361_un1_Y));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I350_un1_Y (.A(N778), .B(N794), 
        .C(N1097), .Y(I350_un1_Y));
    VCC VCC_i (.Y(VCC));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I221_Y (.A(N698), .B(N706), .Y(
        N780));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I14_G0N (.A(\un1_next_sum[14] )
        , .B(sum_14), .Y(N513_0));
    OR2 \preg_RNI1E1L3[12]  (.A(\un1_next_sum_iv_2[12] ), .B(
        \un1_next_sum_iv_1[12] ), .Y(\un1_next_sum[12] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I116_Y (.A(N471), .B(I116_un1_Y), 
        .Y(N666));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I50_Y (.A(\sumreg[32]_net_1 ), 
        .B(\sumreg[33]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N600)
        );
    AND3 inf_abs1_a_2_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(
        \DWACT_FINC_E[4] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I6_G0N (.A(\un1_next_sum[6] ), 
        .B(sum_6), .Y(N489));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I385_Y_1 (.A(N768), .B(N783), .C(
        ADD_40x40_fast_I385_Y_0), .Y(ADD_40x40_fast_I385_Y_1));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I309_Y (.A(N812), .B(N796), .Y(
        N880));
    AO1 next_ireg_3_0_ADD_22x22_fast_I130_Y (.A(
        ADD_22x22_fast_I130_un1_Y_0), .B(N394), .C(
        ADD_22x22_fast_I130_Y_0), .Y(N510));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I383_un1_Y (.A(N880), .B(N745), 
        .C(N848), .Y(I383_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I185_Y (.A(N661), .B(N657), .Y(
        N738));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I448_Y_0 (.A(
        \sumreg[30]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I448_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I107_Y (.A(N487), .B(N484), .Y(
        N657));
    AO1 next_ireg_3_0_ADD_22x22_fast_I129_Y_0 (.A(N384), .B(N377), .C(
        N376), .Y(ADD_22x22_fast_I129_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I228_Y (.A(N713), .B(N706), .C(
        N705), .Y(N787));
    NOR3B \ireg_RNIJBDP[14]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[14]_net_1 ), .Y(\un3_next_sum_m[14] ));
    NOR3 inf_abs1_a_2_I_8 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2]), 
        .Y(N_11_1));
    NOR2B \preg_RNI8RBI_0[14]  (.A(\preg[14]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[14] ));
    XA1B \sumreg_RNO[26]  (.A(N1052), .B(ADD_40x40_fast_I444_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[26] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I454_Y_0 (.A(
        \sumreg[36]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I454_Y_0));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I110_Y (.A(sum_3), .B(sum_2_d0), 
        .C(\un1_next_sum[0] ), .Y(N660));
    XA1B \sumreg_RNO[17]  (.A(N1079), .B(ADD_40x40_fast_I435_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[17] ));
    NOR3B \ireg_RNI6CKH[6]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[6]_net_1 ), .Y(\un3_next_sum_m[6] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I286_un1_Y (.A(N789), .B(N774), 
        .Y(I286_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I359_Y (.A(N880), .B(N745), .C(
        N879), .Y(N1076));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I137_Y (.A(N609), .B(N613), .Y(
        N690));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I129_un1_Y_0 (.A(N377), .B(N385)
        , .Y(ADD_22x22_fast_I129_un1_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I453_Y_0 (.A(
        \sumreg[35]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I453_Y_0));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I48_Y (.A(\sumreg[33]_net_1 ), 
        .B(\sumreg[34]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N598)
        );
    NOR2A inf_abs1_a_2_I_25 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .Y(
        N_5));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I157_Y (.A(N629), .B(N633), .Y(
        N710));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I428_Y_0 (.A(sum_10), .B(
        \un1_next_sum[10] ), .Y(ADD_40x40_fast_I428_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I312_Y (.A(N815), .B(N800), .C(
        N799), .Y(N883));
    DFN1E1C0 \preg[11]  (.D(\p_adj[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[11]_net_1 ));
    XA1B \sumreg_RNO[23]  (.A(N1061), .B(ADD_40x40_fast_I441_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[23] ));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I131_un1_Y (.A(N389), .B(N381), 
        .C(N396), .Y(I131_un1_Y));
    DFN1E1C0 \sumreg[22]  (.D(\next_sum[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_22));
    OR2 next_ireg_3_0_ADD_22x22_fast_I115_Y (.A(I115_un1_Y), .B(N392), 
        .Y(N531));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I5_P0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[5] ), .C(sum_5), .Y(N487));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I20_G0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[20] ), .C(sum_20), .Y(N531_0));
    DFN1E1C0 \ireg[13]  (.D(\next_ireg_3[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[13]_net_1 ));
    XA1B \sumreg_RNO[29]  (.A(N1043), .B(ADD_40x40_fast_I447_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[29] ));
    DFN1E1C0 \p_adj[8]  (.D(\inf_abs1_5[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[8]_net_1 ));
    OR2 \preg_RNIB8ST2[6]  (.A(\un1_next_sum_iv_2[6] ), .B(
        \un1_next_sum_iv_1[6] ), .Y(\un1_next_sum[6] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I61_Y (.A(N330), .B(N334), .Y(
        N369));
    AX1D next_ireg_3_0_ADD_22x22_fast_I177_Y (.A(I124_un1_Y), .B(
        ADD_22x22_fast_I144_Y_2), .C(ADD_22x22_fast_I177_Y_0), .Y(
        \next_ireg_3[23] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I84_Y (.A(N357), .B(N354), .C(
        N353), .Y(N392));
    OR3 \preg_RNIKLGV1[11]  (.A(\un24_next_sum_m[11] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[11] ), .Y(
        \un1_next_sum_iv_2[11] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I240_Y (.A(N725), .B(N718), .C(
        N717), .Y(N799));
    XNOR2 inf_abs1_a_2_I_7 (.A(sr_new[2]), .B(N_12), .Y(
        \inf_abs1_a_2[2] ));
    XNOR2 inf_abs2_a_0_I_17 (.A(integral[12]), .B(N_21), .Y(
        \inf_abs2_a_0[6] ));
    DFN1E1C0 \sumreg[12]  (.D(\next_sum[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_12));
    DFN1E1C0 \ireg[15]  (.D(\next_ireg_3[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[15]_net_1 ));
    XA1B \sumreg_RNO[1]  (.A(N666), .B(ADD_40x40_fast_I419_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[1] ));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I179_Y (.A(\i_adj[19]_net_1 ), 
        .B(\i_adj[21]_net_1 ), .C(N492), .Y(\next_ireg_3[25] ));
    OR3 \preg_RNIF9562[16]  (.A(\un24_next_sum_m[16] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[16] ), .Y(
        \un1_next_sum_iv_2[16] ));
    OR2 \preg_RNI87581[6]  (.A(next_sum_0_sqmuxa_1), .B(
        \un24_next_sum_m[6] ), .Y(\un1_next_sum_iv_0[6] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I97_Y (.A(sum_10), .B(
        \un1_next_sum[10] ), .C(N499), .Y(N647));
    OR2 next_ireg_3_0_ADD_22x22_fast_I8_P0N (.A(\i_adj[8]_net_1 ), .B(
        \i_adj[10]_net_1 ), .Y(N291));
    DFN1E1C0 \sumreg_2[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(sum_2_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I7_P0N (.A(\i_adj[7]_net_1 ), .B(
        \i_adj[9]_net_1 ), .Y(N288));
    NOR3 inf_abs1_a_2_I_18 (.A(sr_new[4]), .B(sr_new[3]), .C(sr_new[5])
        , .Y(\DWACT_FINC_E_0[2] ));
    XNOR2 inf_abs1_a_2_I_26 (.A(sr_new[9]), .B(N_5), .Y(
        \inf_abs1_a_2[9] ));
    
endmodule


module sig_gen_5(
       vd_done,
       n_rst_c,
       clk_c,
       vd_rdy
    );
input  vd_done;
input  n_rst_c;
input  clk_c;
output vd_rdy;

    wire sig_prev_i, sig_prev_net_1, sig_old_i_0, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    NOR2B sig_old_RNIICF1 (.A(sig_old_i_0), .B(sig_prev_net_1), .Y(
        vd_rdy));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(clk_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev (.D(vd_done), .CLK(clk_c), .CLR(n_rst_c), .Q(
        sig_prev_net_1));
    INV sig_old_RNO (.A(sig_prev_net_1), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module spi_stp_12s_1_6_1(
       cur_vd,
       N_29,
       din_5_c,
       n_rst_c,
       sck_fb_c
    );
output [11:0] cur_vd;
input  N_29;
input  din_5_c;
input  n_rst_c;
input  sck_fb_c;

    wire GND, VCC;
    
    DFN1E0C0 \sr[7]  (.D(cur_vd[6]), .CLK(sck_fb_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[7]));
    DFN1E0C0 \sr[5]  (.D(cur_vd[4]), .CLK(sck_fb_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[5]));
    DFN1E0C0 \sr[10]  (.D(cur_vd[9]), .CLK(sck_fb_c), .CLR(n_rst_c), 
        .E(N_29), .Q(cur_vd[10]));
    DFN1E0C0 \sr[8]  (.D(cur_vd[7]), .CLK(sck_fb_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[8]));
    DFN1E0C0 \sr[3]  (.D(cur_vd[2]), .CLK(sck_fb_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[3]));
    DFN1E0C0 \sr[1]  (.D(cur_vd[0]), .CLK(sck_fb_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[1]));
    DFN1E0C0 \sr[2]  (.D(cur_vd[1]), .CLK(sck_fb_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[2]));
    DFN1E0C0 \sr[9]  (.D(cur_vd[8]), .CLK(sck_fb_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[9]));
    VCC VCC_i (.Y(VCC));
    DFN1E0C0 \sr[11]  (.D(cur_vd[10]), .CLK(sck_fb_c), .CLR(n_rst_c), 
        .E(N_29), .Q(cur_vd[11]));
    DFN1E0C0 \sr[0]  (.D(din_5_c), .CLK(sck_fb_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[0]));
    GND GND_i (.Y(GND));
    DFN1E0C0 \sr[6]  (.D(cur_vd[5]), .CLK(sck_fb_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[6]));
    DFN1E0C0 \sr[4]  (.D(cur_vd[3]), .CLK(sck_fb_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[4]));
    
endmodule


module sig_gen_10_4(
       cs_i_1,
       n_rst_c,
       sck_fb_c,
       vd_done
    );
input  cs_i_1;
input  n_rst_c;
input  sck_fb_c;
output vd_done;

    wire sig_prev_i, sig_prev_net_1, sig_old_i_0, GND, VCC;
    
    NOR2B sig_old_RNI8LOE (.A(sig_prev_net_1), .B(sig_old_i_0), .Y(
        vd_done));
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(sck_fb_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev (.D(cs_i_1), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        sig_prev_net_1));
    INV sig_old_RNO (.A(sig_prev_net_1), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module spi_ctl_12s_3_1(
       n_rst_c,
       sck_fb_c,
       N_29,
       cs_i_1,
       cs_i_1_i
    );
input  n_rst_c;
input  sck_fb_c;
output N_29;
output cs_i_1;
output cs_i_1_i;

    wire cnt_m1_0_a2_0, \cnt[14]_net_1 , \cnt[13]_net_1 , 
        cnt_m6_0_a2_6, cnt_m6_0_a2_0, \cnt[3]_net_1 , cnt_m5_0_a2_2, 
        cnt_m6_0_a2_2, \cnt[7]_net_1 , \cnt[8]_net_1 , \cnt[11]_net_1 , 
        \cnt[10]_net_1 , cnt_m7_0_a2_4, \cnt[5]_net_1 , cnt_m7_0_a2_3, 
        \cnt[6]_net_1 , cnt_m7_0_a2_1, \cnt[9]_net_1 , 
        state_tr0_0_a3_12, state_tr0_0_a3_6, state_tr0_0_a3_9, N_103, 
        \cnt[4]_net_1 , state_tr0_0_a3_8, state_tr0_0_a3_3, 
        \cnt[12]_net_1 , state_tr0_0_a3_7, state_tr0_0_a3_2, 
        \cnt[0]_net_1 , \cnt[1]_net_1 , state_tr0_0_a3_1, 
        \cnt[15]_net_1 , vd_stp_en_i_a3_9, vd_stp_en_i_a3_4, N_73, 
        vd_stp_en_i_a3_8, vd_stp_en_i_a3_2, vd_stp_en_i_a3_5, 
        cnt_m6_0_a2_5_6, cnt_m6_0_a2_5_0, cnt_m6_0_a2_5, 
        \cnt[2]_net_1 , cnt_m5_0_a2_3, cnt_m2_0_a2_0, cnt_m5_0_a2_1, 
        cnt_m2_0_a2_2, cnt_m2_0_a2_1, N_74, cnt_N_13_mux, N_33, N_31, 
        cnt_N_7_mux_0_0, cnt_N_3_mux_0, cnt_N_11_mux_2, cnt_N_15_mux, 
        cnt_N_13_mux_0, N_30, \state_RNO_6[0] , N_26, N_24, N_22, N_20, 
        N_97, N_18, N_14, N_12, N_36, \cnt_RNO_1[6]_net_1 , cnt_n10, 
        d_N_3_mux_0, \cnt_RNO_1_2[10] , cnt_n0, N_38, cnt_n15, cnt_n14, 
        cnt_n13, N_72, cnt_n12, cnt_n11, cnt_n9, GND, VCC;
    
    NOR2B \cnt_RNO_2[6]  (.A(\cnt[4]_net_1 ), .B(\cnt[3]_net_1 ), .Y(
        cnt_m2_0_a2_2));
    XA1A \cnt_RNO[8]  (.A(N_36), .B(\cnt[8]_net_1 ), .C(cs_i_1), .Y(
        N_12));
    NOR3C \cnt_RNISP43[4]  (.A(vd_stp_en_i_a3_4), .B(state_tr0_0_a3_3), 
        .C(N_73), .Y(vd_stp_en_i_a3_9));
    NOR3C \cnt_RNO_3[10]  (.A(\cnt[3]_net_1 ), .B(\cnt[5]_net_1 ), .C(
        cs_i_1), .Y(cnt_m7_0_a2_4));
    NOR2B \cnt_RNIFNS[5]  (.A(\cnt[4]_net_1 ), .B(\cnt[5]_net_1 ), .Y(
        cnt_m5_0_a2_2));
    NOR3A \state_RNO_0[0]  (.A(state_tr0_0_a3_3), .B(\cnt[12]_net_1 ), 
        .C(\cnt[9]_net_1 ), .Y(state_tr0_0_a3_8));
    NOR3B \cnt_RNIKNP11[3]  (.A(cnt_m6_0_a2_6), .B(cnt_m6_0_a2_5), .C(
        N_31), .Y(cnt_N_13_mux));
    XA1A \cnt_RNO[2]  (.A(N_30), .B(\cnt[2]_net_1 ), .C(cs_i_1), .Y(
        N_24));
    NOR2B \cnt_RNI7FS_0[1]  (.A(\cnt[1]_net_1 ), .B(\cnt[0]_net_1 ), 
        .Y(cnt_m2_0_a2_0));
    NOR2 \cnt_RNIC5AT[11]  (.A(\cnt[11]_net_1 ), .B(\cnt[13]_net_1 ), 
        .Y(state_tr0_0_a3_1));
    DFN1C0 \cnt[2]  (.D(N_24), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[2]_net_1 ));
    DFN1C0 \cnt[8]  (.D(N_12), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[8]_net_1 ));
    DFN1C0 \cnt[1]  (.D(N_26), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[1]_net_1 ));
    OA1C \cnt_RNO_0[4]  (.A(\cnt[3]_net_1 ), .B(N_31), .C(
        \cnt[4]_net_1 ), .Y(N_97));
    DFN1C0 \cnt[11]  (.D(cnt_n11), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[11]_net_1 ));
    NOR3C \cnt_RNIA743[3]  (.A(cnt_m5_0_a2_2), .B(cnt_m5_0_a2_1), .C(
        cnt_m5_0_a2_3), .Y(cnt_N_11_mux_2));
    NOR3C \cnt_RNO_0[6]  (.A(cnt_m2_0_a2_1), .B(cnt_m2_0_a2_0), .C(
        cnt_m2_0_a2_2), .Y(cnt_N_7_mux_0_0));
    NOR2B \cnt_RNO_1[15]  (.A(\cnt[14]_net_1 ), .B(\cnt[13]_net_1 ), 
        .Y(cnt_m1_0_a2_0));
    XA1A \cnt_RNO[3]  (.A(N_31), .B(\cnt[3]_net_1 ), .C(cs_i_1), .Y(
        N_22));
    OR2B \cnt_RNO_0[13]  (.A(cnt_N_13_mux), .B(\cnt[12]_net_1 ), .Y(
        N_72));
    VCC VCC_i (.Y(VCC));
    XA1 \cnt_RNO[1]  (.A(\cnt[0]_net_1 ), .B(\cnt[1]_net_1 ), .C(
        cs_i_1), .Y(N_26));
    NOR2 \cnt_RNIJRS[6]  (.A(\cnt[7]_net_1 ), .B(\cnt[6]_net_1 ), .Y(
        state_tr0_0_a3_3));
    DFN1C0 \cnt[6]  (.D(\cnt_RNO_1[6]_net_1 ), .CLK(sck_fb_c), .CLR(
        n_rst_c), .Q(\cnt[6]_net_1 ));
    NOR3C \cnt_RNO_0[15]  (.A(cnt_m1_0_a2_0), .B(\cnt[12]_net_1 ), .C(
        cnt_N_13_mux), .Y(cnt_N_3_mux_0));
    NOR3C \cnt_RNIFVCO2[10]  (.A(vd_stp_en_i_a3_2), .B(
        state_tr0_0_a3_1), .C(vd_stp_en_i_a3_5), .Y(vd_stp_en_i_a3_8));
    NOR3A \state_RNO_1[0]  (.A(state_tr0_0_a3_2), .B(\cnt[0]_net_1 ), 
        .C(\cnt[1]_net_1 ), .Y(state_tr0_0_a3_7));
    DFN1C0 \cnt[4]  (.D(N_20), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[4]_net_1 ));
    DFN1C0 \cnt[9]  (.D(cnt_n9), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[9]_net_1 ));
    NOR2A \cnt_RNO[0]  (.A(cs_i_1), .B(\cnt[0]_net_1 ), .Y(cnt_n0));
    NOR2 \cnt_RNIA3AT[10]  (.A(\cnt[10]_net_1 ), .B(\cnt[12]_net_1 ), 
        .Y(vd_stp_en_i_a3_2));
    OR3C \cnt_RNO_0[14]  (.A(\cnt[12]_net_1 ), .B(\cnt[13]_net_1 ), .C(
        cnt_N_13_mux), .Y(N_74));
    AO1B \state_RNIAHR33[0]  (.A(vd_stp_en_i_a3_9), .B(
        vd_stp_en_i_a3_8), .C(cs_i_1), .Y(N_29));
    DFN1C0 \cnt[0]  (.D(cnt_n0), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[0]_net_1 ));
    NOR3B \cnt_RNO[4]  (.A(N_33), .B(cs_i_1), .C(N_97), .Y(N_20));
    NOR3A \state_RNO_4[0]  (.A(state_tr0_0_a3_1), .B(\cnt[14]_net_1 ), 
        .C(\cnt[15]_net_1 ), .Y(state_tr0_0_a3_6));
    NOR2 \cnt_RNIBJS[2]  (.A(\cnt[3]_net_1 ), .B(\cnt[2]_net_1 ), .Y(
        N_103));
    DFN1C0 \state[0]  (.D(\state_RNO_6[0] ), .CLK(sck_fb_c), .CLR(
        n_rst_c), .Q(cs_i_1));
    NOR2B \cnt_RNI92AT[11]  (.A(\cnt[11]_net_1 ), .B(\cnt[10]_net_1 ), 
        .Y(cnt_m6_0_a2_0));
    XA1 \cnt_RNO[6]  (.A(cnt_N_7_mux_0_0), .B(\cnt[6]_net_1 ), .C(
        cs_i_1), .Y(\cnt_RNO_1[6]_net_1 ));
    XA1 \cnt_RNO[15]  (.A(\cnt[15]_net_1 ), .B(cnt_N_3_mux_0), .C(
        cs_i_1), .Y(cnt_n15));
    XA1A \cnt_RNO[9]  (.A(\cnt[9]_net_1 ), .B(N_38), .C(cs_i_1), .Y(
        cnt_n9));
    GND GND_i (.Y(GND));
    NOR2B \cnt_RNO_5[10]  (.A(\cnt[8]_net_1 ), .B(\cnt[9]_net_1 ), .Y(
        cnt_m7_0_a2_1));
    INV \state_RNIVN98[0]  (.A(cs_i_1), .Y(cs_i_1_i));
    DFN1C0 \cnt[13]  (.D(cnt_n13), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[13]_net_1 ));
    NOR3B \state_RNO_5[0]  (.A(\cnt[5]_net_1 ), .B(N_103), .C(
        \cnt[4]_net_1 ), .Y(state_tr0_0_a3_9));
    NOR2B \cnt_RNIDPA1[3]  (.A(\cnt[3]_net_1 ), .B(cnt_m2_0_a2_0), .Y(
        cnt_m5_0_a2_3));
    OR2A \cnt_RNO_0[9]  (.A(\cnt[8]_net_1 ), .B(N_36), .Y(N_38));
    OR2A \cnt_RNICOA1[2]  (.A(\cnt[2]_net_1 ), .B(N_30), .Y(N_31));
    DFN1C0 \cnt[7]  (.D(N_14), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[7]_net_1 ));
    NOR3C \state_RNO_2[0]  (.A(state_tr0_0_a3_6), .B(cs_i_1), .C(
        state_tr0_0_a3_9), .Y(state_tr0_0_a3_12));
    OR3B \cnt_RNIPD72[4]  (.A(\cnt[3]_net_1 ), .B(\cnt[4]_net_1 ), .C(
        N_31), .Y(N_33));
    DFN1C0 \cnt[10]  (.D(cnt_n10), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[10]_net_1 ));
    NOR3C \cnt_RNO_1[11]  (.A(cnt_m6_0_a2_5_0), .B(\cnt[3]_net_1 ), .C(
        cnt_m5_0_a2_2), .Y(cnt_m6_0_a2_5_6));
    XA1A \cnt_RNO[5]  (.A(N_33), .B(\cnt[5]_net_1 ), .C(cs_i_1), .Y(
        N_18));
    NOR3 \cnt_RNIPMOT[15]  (.A(\cnt[14]_net_1 ), .B(\cnt[15]_net_1 ), 
        .C(\cnt[5]_net_1 ), .Y(vd_stp_en_i_a3_5));
    NOR2 \cnt_RNINVS[9]  (.A(\cnt[9]_net_1 ), .B(\cnt[8]_net_1 ), .Y(
        vd_stp_en_i_a3_4));
    OR2B \cnt_RNI7FS[1]  (.A(\cnt[1]_net_1 ), .B(\cnt[0]_net_1 ), .Y(
        N_30));
    NOR3C \cnt_RNIU3LU[3]  (.A(cnt_m6_0_a2_0), .B(\cnt[3]_net_1 ), .C(
        cnt_m5_0_a2_2), .Y(cnt_m6_0_a2_6));
    NOR2B \cnt_RNILTS[7]  (.A(\cnt[7]_net_1 ), .B(\cnt[8]_net_1 ), .Y(
        cnt_m6_0_a2_2));
    NOR2B \cnt_RNIEMS[6]  (.A(\cnt[2]_net_1 ), .B(\cnt[6]_net_1 ), .Y(
        cnt_m5_0_a2_1));
    DFN1C0 \cnt[3]  (.D(N_22), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[3]_net_1 ));
    NOR2B \cnt_RNO_2[11]  (.A(\cnt[10]_net_1 ), .B(\cnt[2]_net_1 ), .Y(
        cnt_m6_0_a2_5_0));
    XA1A \cnt_RNO[14]  (.A(\cnt[14]_net_1 ), .B(N_74), .C(cs_i_1), .Y(
        cnt_n14));
    XNOR2 \cnt_RNO_1[10]  (.A(\cnt[10]_net_1 ), .B(\cnt[4]_net_1 ), .Y(
        \cnt_RNO_1_2[10] ));
    NOR3C \cnt_RNO_4[10]  (.A(\cnt[7]_net_1 ), .B(\cnt[6]_net_1 ), .C(
        cnt_m7_0_a2_1), .Y(cnt_m7_0_a2_3));
    NOR3B \cnt_RNO_0[11]  (.A(cnt_m6_0_a2_5), .B(cnt_m6_0_a2_5_6), .C(
        N_30), .Y(cnt_N_13_mux_0));
    XA1 \cnt_RNO[11]  (.A(\cnt[11]_net_1 ), .B(cnt_N_13_mux_0), .C(
        cs_i_1), .Y(cnt_n11));
    NOR3B \cnt_RNO_2[10]  (.A(cnt_m7_0_a2_4), .B(cnt_m7_0_a2_3), .C(
        N_31), .Y(cnt_N_15_mux));
    OR2A \cnt_RNIIUA1[4]  (.A(\cnt[4]_net_1 ), .B(N_103), .Y(N_73));
    OR3C \state_RNO[0]  (.A(state_tr0_0_a3_8), .B(state_tr0_0_a3_7), 
        .C(state_tr0_0_a3_12), .Y(\state_RNO_6[0] ));
    MX2B \cnt_RNO[10]  (.A(d_N_3_mux_0), .B(\cnt_RNO_1_2[10] ), .S(
        cnt_N_15_mux), .Y(cnt_n10));
    DFN1C0 \cnt[15]  (.D(cnt_n15), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[15]_net_1 ));
    OR2B \cnt_RNIKLI3[7]  (.A(\cnt[7]_net_1 ), .B(cnt_N_11_mux_2), .Y(
        N_36));
    NOR2B \cnt_RNO_1[6]  (.A(\cnt[2]_net_1 ), .B(\cnt[5]_net_1 ), .Y(
        cnt_m2_0_a2_1));
    NOR2B \cnt_RNO_0[10]  (.A(\cnt[10]_net_1 ), .B(cs_i_1), .Y(
        d_N_3_mux_0));
    NOR2 \state_RNO_3[0]  (.A(\cnt[10]_net_1 ), .B(\cnt[8]_net_1 ), .Y(
        state_tr0_0_a3_2));
    NOR3C \cnt_RNIARP1[6]  (.A(\cnt[9]_net_1 ), .B(\cnt[6]_net_1 ), .C(
        cnt_m6_0_a2_2), .Y(cnt_m6_0_a2_5));
    DFN1C0 \cnt[5]  (.D(N_18), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[5]_net_1 ));
    XA1A \cnt_RNO[13]  (.A(\cnt[13]_net_1 ), .B(N_72), .C(cs_i_1), .Y(
        cnt_n13));
    XA1 \cnt_RNO[12]  (.A(\cnt[12]_net_1 ), .B(cnt_N_13_mux), .C(
        cs_i_1), .Y(cnt_n12));
    DFN1C0 \cnt[12]  (.D(cnt_n12), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[12]_net_1 ));
    XA1 \cnt_RNO[7]  (.A(cnt_N_11_mux_2), .B(\cnt[7]_net_1 ), .C(
        cs_i_1), .Y(N_14));
    DFN1C0 \cnt[14]  (.D(cnt_n14), .CLK(sck_fb_c), .CLR(n_rst_c), .Q(
        \cnt[14]_net_1 ));
    
endmodule


module spi_rx_12s_2(
       cur_vd,
       vd_done,
       cs_i_1_i,
       sck_fb_c,
       n_rst_c,
       din_5_c
    );
output [11:0] cur_vd;
output vd_done;
output cs_i_1_i;
input  sck_fb_c;
input  n_rst_c;
input  din_5_c;

    wire N_29, cs_i_1, GND, VCC;
    
    spi_stp_12s_1_6_1 VD_STP (.cur_vd({cur_vd[11], cur_vd[10], 
        cur_vd[9], cur_vd[8], cur_vd[7], cur_vd[6], cur_vd[5], 
        cur_vd[4], cur_vd[3], cur_vd[2], cur_vd[1], cur_vd[0]}), .N_29(
        N_29), .din_5_c(din_5_c), .n_rst_c(n_rst_c), .sck_fb_c(
        sck_fb_c));
    sig_gen_10_4 SPI_RDYSIG (.cs_i_1(cs_i_1), .n_rst_c(n_rst_c), 
        .sck_fb_c(sck_fb_c), .vd_done(vd_done));
    VCC VCC_i (.Y(VCC));
    spi_ctl_12s_3_1 SPICTL (.n_rst_c(n_rst_c), .sck_fb_c(sck_fb_c), 
        .N_29(N_29), .cs_i_1(cs_i_1), .cs_i_1_i(cs_i_1_i));
    GND GND_i (.Y(GND));
    
endmodule


module integral_calc_13s_0_4_2(
       sr_new,
       sr_old,
       sr_new_0_0,
       sr_new_1_0,
       integral,
       integral_i,
       integral_0_0,
       integral_1_0,
       calc_int,
       N_46_1,
       n_rst_c,
       clk_c
    );
input  [12:0] sr_new;
input  [12:0] sr_old;
input  sr_new_0_0;
input  sr_new_1_0;
output [25:6] integral;
output [25:24] integral_i;
output integral_0_0;
output integral_1_0;
input  calc_int;
output N_46_1;
input  n_rst_c;
input  clk_c;

    wire \un1_integ[25] , \un1_next_int_0_iv_0[13] , next_int_1_sqmuxa, 
        next_int_0_sqmuxa_1, N_46_1_0, \state[0]_net_1 , 
        \state[1]_net_1 , N_12, N_10, \DWACT_FINC_E[0] , N_5, 
        \DWACT_FINC_E[4] , N_2, \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , 
        N_12_0, N_10_0, \DWACT_FINC_E_0[0] , N_5_0, 
        \DWACT_FINC_E_0[4] , N_2_0, \DWACT_FINC_E_0[7] , 
        \DWACT_FINC_E_0[6] , ADD_26x26_fast_I255_Y_0, 
        \un1_next_int_0_iv[13] , ADD_26x26_fast_I254_Y_0, 
        ADD_26x26_fast_I253_Y_0, ADD_26x26_fast_I252_Y_0, 
        ADD_26x26_fast_I249_Y_0, ADD_26x26_fast_I246_Y_0, 
        ADD_26x26_fast_I247_Y_0, ADD_26x26_fast_I204_Y_3, N502, N517, 
        ADD_26x26_fast_I204_Y_2, N398, ADD_26x26_fast_I204_Y_0, N455, 
        ADD_26x26_fast_I205_Y_3, N504, N519, ADD_26x26_fast_I205_Y_2, 
        N400, ADD_26x26_fast_I205_Y_0, N457, ADD_26x26_fast_I248_Y_0, 
        ADD_26x26_fast_I250_Y_0, ADD_26x26_fast_I251_Y_0, 
        ADD_26x26_fast_I206_Y_2, ADD_26x26_fast_I206_un1_Y_0, N522, 
        ADD_26x26_fast_I206_Y_1, I80_un1_Y, N459, 
        ADD_26x26_fast_I245_Y_0, ADD_26x26_fast_I207_Y_2, 
        ADD_26x26_fast_I207_un1_Y_0, N524, ADD_26x26_fast_I207_Y_1, 
        N404, N461, ADD_26x26_fast_I210_Y_1, N514, N529, 
        ADD_26x26_fast_I210_Y_0, N467, N460, ADD_26x26_fast_I212_Y_0, 
        N533, N518, ADD_26x26_fast_I213_Y_0, N535, N520, 
        ADD_26x26_fast_I242_Y_0, \un2_next_int_m[12] , 
        \un1_next_int_iv_0[12] , ADD_26x26_fast_I244_Y_0, 
        ADD_26x26_fast_I241_Y_0, \un1_next_int[11] , 
        ADD_26x26_fast_I243_Y_0, ADD_26x26_fast_I211_Y_0, N469, N462, 
        ADD_26x26_fast_I208_Y_1, ADD_26x26_fast_I208_un1_Y_0, N526, 
        ADD_26x26_fast_I208_Y_0, N463, ADD_26x26_fast_I209_Y_1, 
        ADD_26x26_fast_I209_un1_Y_0, N528, ADD_26x26_fast_I209_Y_0, 
        N465, N458, ADD_26x26_fast_I204_un1_Y_0, 
        ADD_26x26_fast_I205_un1_Y_0, ADD_26x26_fast_I239_Y_0, 
        \un2_next_int_m[9] , \un1_next_int_iv_1[9] , 
        ADD_26x26_fast_I240_Y_0, \un1_next_int[10] , 
        ADD_26x26_fast_I238_Y_0, \un1_next_int[8] , 
        ADD_26x26_fast_I211_Y_1_0, N470, ADD_26x26_fast_I213_un1_Y_0, 
        N482, N490, \un1_next_int[0] , N483, I160_un1_Y, N506, N485, 
        I161_un1_Y, N508, N487, I162_un1_Y, N510, N489, I163_un1_Y, 
        N512, ADD_26x26_fast_I237_Y_0, \un1_next_int[7] , 
        ADD_26x26_fast_I235_Y_0, \integ[5]_net_1 , \un1_next_int[5] , 
        ADD_26x26_fast_I236_Y_0, \un1_next_int[6] , 
        ADD_26x26_fast_I234_Y_0, \integ[4]_net_1 , \un1_next_int[4] , 
        ADD_26x26_fast_I232_Y_0, \integ[2]_net_1 , \un1_next_int[2] , 
        ADD_26x26_fast_I127_Y_0, ADD_26x26_fast_I125_Y_0, 
        ADD_26x26_fast_I231_Y_0, \integ[1]_net_1 , \un1_next_int[1] , 
        \un1_next_int_iv_0[11] , \inf_abs1[11]_net_1 , 
        \un1_next_int_iv_0[10] , \inf_abs1[10]_net_1 , 
        \inf_abs1_a_1[12] , \un1_next_int_iv_1[4] , 
        \un1_next_int_iv_0[4] , \inf_abs0_m[4] , \inf_abs1[4]_net_1 , 
        \un1_next_int_iv_0[8] , \inf_abs1[8]_net_1 , 
        \un1_next_int_iv_0[6] , \inf_abs1[6]_net_1 , 
        ADD_26x26_fast_I230_Y_0, \integ[0]_net_1 , N_3, 
        \inf_abs0_m[9] , \un18_next_int_m[9] , \inf_abs1_m[9] , 
        \un1_next_int_iv_1[0] , \un1_next_int_iv_0[0] , 
        \inf_abs0_m[0] , \un18_next_int_m[0] , \inf_abs1_m[0] , 
        \un1_next_int_iv_1[5] , \inf_abs0_m[5] , \un18_next_int_m[5] , 
        \inf_abs1_m[5] , \un1_next_int_iv_1[7] , \inf_abs0_m[7] , 
        \un18_next_int_m[7] , \inf_abs1_m[7] , \un1_next_int_iv_1[1] , 
        \un1_next_int_iv_0[1] , \inf_abs0_m[1] , \un18_next_int_m[1] , 
        \inf_abs1_m[1] , \un1_next_int_iv_1[3] , \inf_abs1_m[3] , 
        \un18_next_int_m[3] , \inf_abs0_m[3] , \un1_next_int_iv_1[2] , 
        \inf_abs1_m[2] , \un18_next_int_m[2] , \inf_abs0_m[2] , 
        ADD_26x26_fast_I211_Y_1, ADD_26x26_fast_I211_un1_Y_0, N531, 
        N399, N456, I204_un1_Y, I194_un1_Y, \un2_next_int_m[5] , 
        \un2_next_int_m[1] , \un2_next_int_m[0] , \un1_integ[5] , 
        \un1_integ[9] , \un2_next_int_m[7] , \un1_next_int[3] , 
        \un2_next_int_m[3] , \un2_next_int_m[2] , \un1_integ[20] , 
        I178_un1_Y, \un1_integ[23] , I172_un1_Y, \un1_integ[13] , N525, 
        I190_un1_Y, \un1_integ[6] , \un1_integ[12] , N527, I191_un1_Y, 
        \un1_integ[14] , N523, I189_un1_Y, \un1_integ[16] , I213_un1_Y, 
        \un1_integ[17] , I212_un1_Y, \un1_integ[24] , I205_un1_Y, 
        \un1_integ[0] , \un1_integ[3] , \integ[3]_net_1 , N491, 
        \un1_integ[7] , \un1_integ[15] , N521, I188_un1_Y, 
        \un1_integ[18] , \un1_integ[19] , I210_un1_Y, \un1_integ[21] , 
        I176_un1_Y, \un1_integ[2] , N493, \un1_integ[10] , I193_un1_Y, 
        \un1_integ[22] , I174_un1_Y, \un1_integ[11] , I192_un1_Y, 
        \un1_integ[8] , I195_un1_Y, \un1_integ[4] , \un1_integ[1] , 
        N442, \un2_next_int_m[4] , \inf_abs0_m[6] , 
        \un2_next_int_m[6] , \inf_abs0_m[8] , \un2_next_int_m[8] , 
        \inf_abs0_m[10] , \un2_next_int_m[10] , \inf_abs0_m[11] , 
        \un2_next_int_m[11] , N530, N403, N534, N405, N401, N478, N486, 
        N474, N481, N480, N479, N430, N427, N426, N338, N339, N488, 
        N439, N321, I150_un1_Y, N473, N424, N421, N420, N347, N351, 
        N350, N348, N425, N345, I146_un1_Y, N417, N416, N353, N354, 
        N477, N429, N466, N413, N412, N419, N423, N464, N411, N415, 
        N471, N440, N437, N436, N327, N441, N318, N433, I110_un1_Y, 
        N428, I60_un1_Y, N335, N432, N409, N408, I74_un1_Y, N317, N422, 
        N418, N475, N476, I144_un1_Y, I148_un1_Y, N484, N414, N438, 
        N320, N323, N344, I56_un1_Y, I106_un1_Y, I121_un1_Y, 
        \inf_abs0[4]_net_1 , \inf_abs0[6]_net_1 , \inf_abs0[8]_net_1 , 
        \inf_abs0[10]_net_1 , \inf_abs0[11]_net_1 , \inf_abs0_a_0[12] , 
        \state_RNO_6[1] , \inf_abs0_a_0[4] , \inf_abs0_a_0[6] , 
        \inf_abs0_a_0[8] , \inf_abs0_a_0[10] , \inf_abs0_a_0[11] , 
        \inf_abs1_a_1[4] , \inf_abs1_a_1[6] , \inf_abs1_a_1[8] , 
        \inf_abs1_a_1[10] , \inf_abs1_a_1[11] , \state_RNO_5[0] , N406, 
        N410, N407, \inf_abs1_a_1[2] , \inf_abs0_a_0[2] , 
        \inf_abs1_a_1[7] , \inf_abs0_a_0[7] , \inf_abs1_a_1[3] , 
        \inf_abs0_a_0[3] , N326, N435, N330, N333, N434, N329, 
        I64_un1_Y, N332, \inf_abs1_a_1[1] , \inf_abs0_a_0[1] , 
        \inf_abs1_a_1[9] , \inf_abs0_a_0[9] , \inf_abs1_a_1[5] , 
        \inf_abs0_a_0[5] , N431, N_3_0, \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[5] , N_4, \DWACT_FINC_E[3] , N_6, N_7, N_8, 
        \DWACT_FINC_E[1] , N_9, N_11, N_3_1, \DWACT_FINC_E_0[2] , 
        \DWACT_FINC_E_0[5] , N_4_0, \DWACT_FINC_E_0[3] , N_6_0, N_7_0, 
        N_8_0, \DWACT_FINC_E_0[1] , N_9_0, N_11_0, GND, VCC;
    
    OR2 un1_integ_0_0_ADD_26x26_fast_I56_Y (.A(I56_un1_Y), .B(N344), 
        .Y(N424));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I148_un1_Y (.A(N419), .B(N423), 
        .C(N479), .Y(I148_un1_Y));
    NOR2 inf_abs1_a_1_I_15 (.A(sr_old[3]), .B(sr_old[4]), .Y(
        \DWACT_FINC_E[1] ));
    XNOR2 inf_abs1_a_1_I_23 (.A(sr_old[8]), .B(N_6), .Y(
        \inf_abs1_a_1[8] ));
    DFN1C0 \state[0]  (.D(\state_RNO_5[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[0]_net_1 ));
    XNOR2 inf_abs1_a_1_I_17 (.A(sr_old[6]), .B(N_8), .Y(
        \inf_abs1_a_1[6] ));
    NOR2B \state_RNIE5RA3[1]  (.A(\inf_abs1_a_1[5] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[5] ));
    DFN1E0C0 \integ[13]  (.D(\un1_integ[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[13]));
    DFN1E0C0 \integ[24]  (.D(\un1_integ[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[24]));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I245_Y_0 (.A(integral[15]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I245_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I61_Y (.A(integral[6]), .B(
        \un1_next_int[6] ), .C(N339), .Y(N429));
    OR2 un1_integ_0_0_ADD_26x26_fast_I7_P0N (.A(\un1_next_int[7] ), .B(
        integral[7]), .Y(N339));
    NOR3B inf_abs0_a_0_I_19 (.A(\DWACT_FINC_E_0[2] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[6]), .Y(N_7_0));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I248_Y_0 (.A(integral[18]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I248_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I172_un1_Y (.A(N506), .B(N521), 
        .Y(I172_un1_Y));
    OR2 \state_RNI74CD7[0]  (.A(\un1_next_int_iv_1[5] ), .B(
        \un2_next_int_m[5] ), .Y(\un1_next_int[5] ));
    NOR3B inf_abs0_a_0_I_16 (.A(\DWACT_FINC_E_0[1] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[5]), .Y(N_8_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I41_Y (.A(integral[17]), .B(
        integral[16]), .C(\un1_next_int_0_iv_0[13] ), .Y(N409));
    OA1 un1_integ_0_0_ADD_26x26_fast_I204_un1_Y (.A(N533), .B(
        I194_un1_Y), .C(ADD_26x26_fast_I204_un1_Y_0), .Y(I204_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I86_Y (.A(N408), .B(N404), .Y(
        N457));
    NOR3A \state_RNIH8P91[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .C(sr_old[7]), .Y(\un18_next_int_m[7] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I98_Y (.A(N420), .B(N417), .C(
        N416), .Y(N469));
    OR3 \state_RNIVIRAB[0]  (.A(\inf_abs0_m[8] ), .B(
        \un1_next_int_iv_0[8] ), .C(\un2_next_int_m[8] ), .Y(
        \un1_next_int[8] ));
    OR2 \state_RNINJ2M8[0]  (.A(\un1_next_int_iv_1[7] ), .B(
        \un2_next_int_m[7] ), .Y(\un1_next_int[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I176_un1_Y (.A(N510), .B(N525), 
        .Y(I176_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I205_un1_Y_0 (.A(N504), .B(N520)
        , .Y(ADD_26x26_fast_I205_un1_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I150_un1_Y (.A(N481), .B(N474), 
        .Y(I150_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I51_Y (.A(N354), .B(N351), .Y(
        N419));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y (.A(
        ADD_26x26_fast_I230_Y_0), .B(\un1_next_int[0] ), .Y(
        \un1_integ[0] ));
    NOR2B \state_RNIJCB03[0]  (.A(\inf_abs0[11]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[11] ));
    NOR2B inf_abs1_a_1_I_34 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .Y(N_2_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I144_un1_Y (.A(N419), .B(N415), 
        .C(N475), .Y(I144_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I253_Y (.A(I172_un1_Y), .B(
        ADD_26x26_fast_I206_Y_2), .C(ADD_26x26_fast_I253_Y_0), .Y(
        \un1_integ[23] ));
    DFN1E0C0 \integ[21]  (.D(\un1_integ[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[21]));
    XNOR2 inf_abs1_a_1_I_7 (.A(sr_old[2]), .B(N_12_0), .Y(
        \inf_abs1_a_1[2] ));
    DFN1E0C0 \integ_1[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral_1_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I190_un1_Y (.A(N487), .B(
        I162_un1_Y), .C(N526), .Y(I190_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I146_Y (.A(I146_un1_Y), .B(N469), 
        .Y(N523));
    AO1 un1_integ_0_0_ADD_26x26_fast_I142_Y (.A(N473), .B(N466), .C(
        N465), .Y(N519));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I244_Y_0 (.A(integral[14]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I244_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I231_Y (.A(
        ADD_26x26_fast_I231_Y_0), .B(N442), .Y(\un1_integ[1] ));
    NOR2B \state_RNIPMOS[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), .Y(
        next_int_0_sqmuxa_1));
    AND3 inf_abs1_a_1_I_24 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E_0[4] ));
    XNOR2 inf_abs1_a_1_I_32 (.A(sr_old[11]), .B(N_3_0), .Y(
        \inf_abs1_a_1[11] ));
    DFN1E0C0 \integ[15]  (.D(\un1_integ[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[15]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I213_un1_Y (.A(
        ADD_26x26_fast_I213_un1_Y_0), .B(N520), .Y(I213_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I103_Y (.A(N425), .B(N421), .Y(
        N474));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I125_Y (.A(N399), .B(
        ADD_26x26_fast_I125_Y_0), .C(N456), .Y(N502));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_1 (.A(
        ADD_26x26_fast_I209_un1_Y_0), .B(N528), .C(
        ADD_26x26_fast_I209_Y_0), .Y(ADD_26x26_fast_I209_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I94_Y (.A(N416), .B(N413), .C(
        N412), .Y(N465));
    NOR2 inf_abs0_a_0_I_6 (.A(sr_new[0]), .B(sr_new[1]), .Y(N_12));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I151_Y (.A(N482), .B(N474), .Y(
        N528));
    AND3 inf_abs1_a_1_I_22 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_6));
    OR2 un1_integ_0_0_ADD_26x26_fast_I74_Y (.A(I74_un1_Y), .B(N317), 
        .Y(N442));
    AX1D un1_integ_0_0_ADD_26x26_fast_I238_Y (.A(N535), .B(I195_un1_Y), 
        .C(ADD_26x26_fast_I238_Y_0), .Y(\un1_integ[8] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I121_Y (.A(I121_un1_Y), .B(N440), 
        .Y(N493));
    OR3 \state_RNIC5676[1]  (.A(\inf_abs0_m[7] ), .B(
        \un18_next_int_m[7] ), .C(\inf_abs1_m[7] ), .Y(
        \un1_next_int_iv_1[7] ));
    NOR3 inf_abs0_a_0_I_10 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2])
        , .Y(\DWACT_FINC_E[0] ));
    NOR2 \state_RNI94SU_0[0]  (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(N_46_1_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I5_P0N (.A(\un1_next_int[5] ), .B(
        \integ[5]_net_1 ), .Y(N333));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I236_Y_0 (.A(integral[6]), .B(
        \un1_next_int[6] ), .Y(ADD_26x26_fast_I236_Y_0));
    NOR3B \state_RNIBESE2[0]  (.A(sr_new_1_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[7] ), .Y(\un2_next_int_m[7] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I246_Y (.A(I213_un1_Y), .B(
        ADD_26x26_fast_I213_Y_0), .C(ADD_26x26_fast_I246_Y_0), .Y(
        \un1_integ[16] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I252_Y_0 (.A(integral[22]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I252_Y_0));
    MX2 \inf_abs0[6]  (.A(sr_new[6]), .B(\inf_abs0_a_0[6] ), .S(
        sr_new_1_0), .Y(\inf_abs0[6]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I39_Y (.A(integral[17]), .B(
        integral[18]), .C(\un1_next_int_0_iv_0[13] ), .Y(N407));
    OA1B un1_integ_0_0_ADD_26x26_fast_I32_Y (.A(integral[21]), .B(
        integral[20]), .C(\un1_next_int_0_iv_0[13] ), .Y(N400));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I194_un1_Y (.A(N534), .B(N442), 
        .Y(I194_un1_Y));
    NOR3B \state_RNIL0IH1[0]  (.A(sr_new_1_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[3] ), .Y(\un2_next_int_m[3] ));
    NOR2A inf_abs0_a_0_I_11 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .Y(
        N_10));
    AO1B un1_integ_0_0_ADD_26x26_fast_I125_Y_0 (.A(integral[23]), .B(
        integral[24]), .C(\un1_next_int_0_iv[13] ), .Y(
        ADD_26x26_fast_I125_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I211_Y_1_0 (.A(N462), .B(N470), 
        .Y(ADD_26x26_fast_I211_Y_1_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I100_Y (.A(N422), .B(N419), .C(
        N418), .Y(N471));
    OR3 un1_integ_0_0_ADD_26x26_fast_I12_P0N (.A(\un2_next_int_m[12] ), 
        .B(\un1_next_int_iv_0[12] ), .C(integral[12]), .Y(N354));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I10_G0N (.A(\un1_next_int[10] ), 
        .B(integral[10]), .Y(N347));
    DFN1E0C0 \integ[12]  (.D(\un1_integ[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[12]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I109_Y (.A(N431), .B(N427), .Y(
        N480));
    XNOR2 inf_abs1_a_1_I_35 (.A(sr_old[12]), .B(N_2_0), .Y(
        \inf_abs1_a_1[12] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I205_Y_0 (.A(integral[22]), .B(
        integral[23]), .C(\un1_next_int_0_iv[13] ), .Y(
        ADD_26x26_fast_I205_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I115_Y (.A(N433), .B(N437), .Y(
        N486));
    NOR3B \state_RNI7HIR_0[0]  (.A(\state[0]_net_1 ), .B(sr_new[0]), 
        .C(sr_new_1_0), .Y(\inf_abs0_m[0] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I12_G0N (.A(\un2_next_int_m[12] ), 
        .B(\un1_next_int_iv_0[12] ), .C(integral[12]), .Y(N353));
    NOR3B \state_RNI2C7V2[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[11]_net_1 ), .Y(\un2_next_int_m[11] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I208_Y_0 (.A(N455), .B(N463), .Y(
        ADD_26x26_fast_I208_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I111_Y (.A(N433), .B(N429), .Y(
        N482));
    NOR2A inf_abs1_a_1_I_25 (.A(\DWACT_FINC_E_0[4] ), .B(sr_old[8]), 
        .Y(N_5_0));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I250_Y_0 (.A(integral[20]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I250_Y_0));
    NOR3A inf_abs1_a_1_I_27 (.A(\DWACT_FINC_E_0[4] ), .B(sr_old[8]), 
        .C(sr_old[9]), .Y(N_4));
    NOR3B \state_RNI9FJU2[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[12] ), .Y(\un2_next_int_m[12] ));
    DFN1E0C0 \integ[10]  (.D(\un1_integ[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[10]));
    NOR2B \state_RNIMO9V2_0[0]  (.A(\inf_abs0[8]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[8] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I188_un1_Y (.A(N483), .B(
        I160_un1_Y), .C(N522), .Y(I188_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I6_G0N (.A(\un1_next_int[6] ), 
        .B(integral[6]), .Y(N335));
    MX2 \inf_abs1[10]  (.A(sr_old[10]), .B(\inf_abs1_a_1[10] ), .S(
        sr_old[12]), .Y(\inf_abs1[10]_net_1 ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I249_Y (.A(I210_un1_Y), .B(
        ADD_26x26_fast_I210_Y_1), .C(ADD_26x26_fast_I249_Y_0), .Y(
        \un1_integ[19] ));
    GND GND_i (.Y(GND));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I146_un1_Y (.A(N477), .B(N470), 
        .Y(I146_un1_Y));
    NOR2B \state_RNIOEGO[0]  (.A(sr_new[1]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[1] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I246_Y_0 (.A(integral[16]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I246_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I1_G0N (.A(\un1_next_int[1] ), 
        .B(\integ[1]_net_1 ), .Y(N320));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I107_Y (.A(N425), .B(N429), .Y(
        N478));
    NOR3B \state_RNI00T21[0]  (.A(sr_new_1_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[1] ), .Y(\un2_next_int_m[1] ));
    XNOR2 inf_abs1_a_1_I_9 (.A(sr_old[3]), .B(N_11), .Y(
        \inf_abs1_a_1[3] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I38_Y (.A(integral[17]), .B(
        integral[18]), .C(\un1_next_int_0_iv_0[13] ), .Y(N406));
    OA1 un1_integ_0_0_ADD_26x26_fast_I209_un1_Y_0 (.A(N489), .B(
        I163_un1_Y), .C(N512), .Y(ADD_26x26_fast_I209_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_3 (.A(N504), .B(N519), .C(
        ADD_26x26_fast_I205_Y_2), .Y(ADD_26x26_fast_I205_Y_3));
    AX1D un1_integ_0_0_ADD_26x26_fast_I255_Y (.A(I204_un1_Y), .B(
        ADD_26x26_fast_I204_Y_3), .C(ADD_26x26_fast_I255_Y_0), .Y(
        \un1_integ[25] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I204_Y_0 (.A(integral[24]), .B(
        integral[23]), .C(\un1_next_int_0_iv_0[13] ), .Y(
        ADD_26x26_fast_I204_Y_0));
    MX2 \inf_abs0[4]  (.A(sr_new[4]), .B(\inf_abs0_a_0[4] ), .S(
        sr_new_0_0), .Y(\inf_abs0[4]_net_1 ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I243_Y (.A(N525), .B(I190_un1_Y), 
        .C(ADD_26x26_fast_I243_Y_0), .Y(\un1_integ[13] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I231_Y_0 (.A(\integ[1]_net_1 ), 
        .B(\un1_next_int[1] ), .Y(ADD_26x26_fast_I231_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I69_Y (.A(\integ[2]_net_1 ), .B(
        \un1_next_int[2] ), .C(N327), .Y(N437));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I62_Y (.A(N332), .B(integral[6]), 
        .C(\un1_next_int[6] ), .Y(N430));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I193_un1_Y (.A(N478), .B(N486), 
        .C(N493), .Y(I193_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I153_Y (.A(N484), .B(N476), .Y(
        N530));
    OR3 \state_RNIPU4D5[1]  (.A(\inf_abs0_m[5] ), .B(
        \un18_next_int_m[5] ), .C(\inf_abs1_m[5] ), .Y(
        \un1_next_int_iv_1[5] ));
    NOR2B \state_RNIQGGO[0]  (.A(sr_new[3]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[3] ));
    XNOR2 inf_abs0_a_0_I_7 (.A(sr_new[2]), .B(N_12), .Y(
        \inf_abs0_a_0[2] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I7_G0N (.A(\un1_next_int[7] ), 
        .B(integral[7]), .Y(N338));
    OA1A un1_integ_0_0_ADD_26x26_fast_I49_Y (.A(
        \un1_next_int_0_iv[13] ), .B(integral[13]), .C(N354), .Y(N417));
    OA1B un1_integ_0_0_ADD_26x26_fast_I42_Y (.A(integral[16]), .B(
        integral[15]), .C(\un1_next_int_0_iv_0[13] ), .Y(N410));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I145_Y (.A(N419), .B(N415), .C(
        N476), .Y(N522));
    NOR2A \state_RNIVV5H[0]  (.A(\state[0]_net_1 ), .B(sr_new[12]), .Y(
        next_int_1_sqmuxa));
    MX2 \inf_abs1[4]  (.A(sr_old[4]), .B(\inf_abs1_a_1[4] ), .S(
        sr_old[12]), .Y(\inf_abs1[4]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I10_P0N (.A(\un1_next_int[10] ), 
        .B(integral[10]), .Y(N348));
    OR2 un1_integ_0_0_ADD_26x26_fast_I1_P0N (.A(\un1_next_int[1] ), .B(
        \integ[1]_net_1 ), .Y(N321));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I192_un1_Y (.A(N530), .B(N491), 
        .Y(I192_un1_Y));
    NOR3A inf_abs0_a_0_I_13 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .C(
        sr_new[4]), .Y(N_9_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I141_Y (.A(N419), .B(N423), .C(
        N464), .Y(N518));
    OA1A \state_RNIP7T66[1]  (.A(sr_old[12]), .B(\inf_abs1_a_1[12] ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[12] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I93_Y (.A(N411), .B(N415), .Y(
        N464));
    AO1B un1_integ_0_0_ADD_26x26_fast_I37_Y (.A(integral[19]), .B(
        integral[18]), .C(\un1_next_int_0_iv_0[13] ), .Y(N405));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I0_G0N (.A(N_3), .B(
        \integ[0]_net_1 ), .Y(N317));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I73_Y (.A(N318), .B(N321), .Y(
        N441));
    OA1 un1_integ_0_0_ADD_26x26_fast_I59_Y (.A(integral[8]), .B(
        \un1_next_int[8] ), .C(N339), .Y(N427));
    AO1 un1_integ_0_0_ADD_26x26_fast_I52_Y (.A(N347), .B(N351), .C(
        N350), .Y(N420));
    NOR2A \state_RNO[1]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 ), 
        .Y(\state_RNO_6[1] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I34_Y (.A(integral[20]), .B(
        integral[19]), .C(\un1_next_int_0_iv_0[13] ), .Y(I80_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I236_Y (.A(N485), .B(I161_un1_Y), 
        .C(ADD_26x26_fast_I236_Y_0), .Y(\un1_integ[6] ));
    NOR2B \state_RNIT7S44[1]  (.A(\inf_abs1_a_1[7] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[7] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I150_Y (.A(I150_un1_Y), .B(N473), 
        .Y(N527));
    NOR2B \state_RNI8EJU2[0]  (.A(\inf_abs0[10]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[10] ));
    DFN1E0C0 \integ[0]  (.D(\un1_integ[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(\integ[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I120_Y (.A(N439), .B(N442), .C(
        N438), .Y(N491));
    AO1 un1_integ_0_0_ADD_26x26_fast_I104_Y (.A(N426), .B(N423), .C(
        N422), .Y(N475));
    VCC VCC_i (.Y(VCC));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I129_Y (.A(N399), .B(N403), .C(
        N460), .Y(N506));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I113_Y (.A(N431), .B(N435), .Y(
        N484));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I241_Y_0 (.A(integral[11]), .B(
        \un1_next_int[11] ), .Y(ADD_26x26_fast_I241_Y_0));
    XNOR2 inf_abs0_a_0_I_28 (.A(sr_new[10]), .B(N_4_0), .Y(
        \inf_abs0_a_0[10] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I89_Y (.A(N407), .B(N411), .Y(
        N460));
    AO1 un1_integ_0_0_ADD_26x26_fast_I68_Y (.A(N323), .B(N327), .C(
        N326), .Y(N436));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_0 (.A(N469), .B(N462), .C(
        N461), .Y(ADD_26x26_fast_I211_Y_0));
    DFN1E0C0 \integ[4]  (.D(\un1_integ[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(\integ[4]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I108_Y (.A(N430), .B(N427), .C(
        N426), .Y(N479));
    NOR2B \state_RNINUOT1[0]  (.A(\inf_abs0[4]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[4] ));
    NOR3 inf_abs1_a_1_I_18 (.A(sr_old[3]), .B(sr_old[5]), .C(sr_old[4])
        , .Y(\DWACT_FINC_E[2] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I3_G0N (.A(\un1_next_int[3] ), 
        .B(\integ[3]_net_1 ), .Y(N326));
    AO13 un1_integ_0_0_ADD_26x26_fast_I48_Y (.A(integral[13]), .B(N353)
        , .C(\un1_next_int_0_iv[13] ), .Y(N416));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I195_un1_Y (.A(N482), .B(N490), 
        .C(\un1_next_int[0] ), .Y(I195_un1_Y));
    DFN1E0C0 \integ[3]  (.D(\un1_integ[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(\integ[3]_net_1 ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I252_Y (.A(I174_un1_Y), .B(
        ADD_26x26_fast_I207_Y_2), .C(ADD_26x26_fast_I252_Y_0), .Y(
        \un1_integ[22] ));
    NOR3B \state_RNIMO9V2[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[8]_net_1 ), .Y(\un2_next_int_m[8] ));
    NOR2B \state_RNISIGO[0]  (.A(sr_new[5]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[5] ));
    DFN1E0C0 \integ[6]  (.D(\un1_integ[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(integral[6]));
    XNOR2 inf_abs0_a_0_I_14 (.A(sr_new[5]), .B(N_9_0), .Y(
        \inf_abs0_a_0[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_1 (.A(N514), .B(N529), .C(
        ADD_26x26_fast_I210_Y_0), .Y(ADD_26x26_fast_I210_Y_1));
    AND3 inf_abs0_a_0_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[5] ), .Y(
        \DWACT_FINC_E[6] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y (.A(N533), .B(I194_un1_Y), 
        .C(ADD_26x26_fast_I239_Y_0), .Y(\un1_integ[9] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I106_un1_Y (.A(N428), .B(N425), 
        .Y(I106_un1_Y));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I58_Y (.A(N338), .B(integral[8]), 
        .C(\un1_next_int[8] ), .Y(N426));
    OR3 \state_RNIKC364[1]  (.A(\inf_abs1_m[2] ), .B(
        \un18_next_int_m[2] ), .C(\inf_abs0_m[2] ), .Y(
        \un1_next_int_iv_1[2] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I67_Y (.A(N330), .B(N327), .Y(
        N435));
    NOR3B \state_RNIQF7A1[0]  (.A(sr_new_1_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[2] ), .Y(\un2_next_int_m[2] ));
    XNOR2 inf_abs0_a_0_I_12 (.A(sr_new[4]), .B(N_10), .Y(
        \inf_abs0_a_0[4] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I253_Y_0 (.A(integral[23]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I253_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I157_Y (.A(N488), .B(N480), .Y(
        N534));
    OR2 un1_integ_0_0_ADD_26x26_fast_I64_Y (.A(I64_un1_Y), .B(N332), 
        .Y(N432));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I204_un1_Y_0 (.A(N502), .B(N518)
        , .Y(ADD_26x26_fast_I204_un1_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I212_un1_Y (.A(N534), .B(N442), 
        .C(N518), .Y(I212_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I127_Y (.A(N401), .B(
        ADD_26x26_fast_I127_Y_0), .C(N458), .Y(N504));
    OR2 un1_integ_0_0_ADD_26x26_fast_I110_Y (.A(I110_un1_Y), .B(N428), 
        .Y(N481));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I211_un1_Y_0 (.A(N478), .B(N486)
        , .C(N493), .Y(ADD_26x26_fast_I211_un1_Y_0));
    OR2 \state_RNIESAG5[0]  (.A(\un1_next_int_iv_1[2] ), .B(
        \un2_next_int_m[2] ), .Y(\un1_next_int[2] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I90_Y (.A(N412), .B(N408), .Y(
        N461));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I233_Y (.A(\un1_next_int[3] ), 
        .B(\integ[3]_net_1 ), .C(N491), .Y(\un1_integ[3] ));
    NOR3A inf_abs0_a_0_I_31 (.A(\DWACT_FINC_E[6] ), .B(sr_new[9]), .C(
        sr_new[10]), .Y(N_3_1));
    AO1B un1_integ_0_0_ADD_26x26_fast_I47_Y (.A(integral[13]), .B(
        integral[14]), .C(\un1_next_int_0_iv_0[13] ), .Y(N415));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I119_Y (.A(N441), .B(N437), .Y(
        N490));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I70_Y (.A(N320), .B(
        \integ[2]_net_1 ), .C(\un1_next_int[2] ), .Y(N438));
    DFN1E0C0 \integ[5]  (.D(\un1_integ[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(\integ[5]_net_1 ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I44_Y (.A(integral[14]), .B(
        integral[15]), .C(\un1_next_int_0_iv_0[13] ), .Y(N412));
    AX1D un1_integ_0_0_ADD_26x26_fast_I245_Y (.A(N521), .B(I188_un1_Y), 
        .C(ADD_26x26_fast_I245_Y_0), .Y(\un1_integ[15] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I95_Y (.A(N413), .B(N417), .Y(
        N466));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y_0 (.A(\un2_next_int_m[9] )
        , .B(\un1_next_int_iv_1[9] ), .C(integral[9]), .Y(
        ADD_26x26_fast_I239_Y_0));
    DFN1E0C0 \integ[2]  (.D(\un1_integ[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(\integ[2]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I135_Y (.A(N458), .B(N466), .Y(
        N512));
    OR2 un1_integ_0_0_ADD_26x26_fast_I88_Y (.A(N406), .B(N410), .Y(
        N459));
    AX1D un1_integ_0_0_ADD_26x26_fast_I247_Y (.A(I212_un1_Y), .B(
        ADD_26x26_fast_I212_Y_0), .C(ADD_26x26_fast_I247_Y_0), .Y(
        \un1_integ[17] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I237_Y_0 (.A(integral[7]), .B(
        \un1_next_int[7] ), .Y(ADD_26x26_fast_I237_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I143_Y (.A(N466), .B(N474), .Y(
        N520));
    NOR2B \state_RNISCPM1[1]  (.A(\inf_abs1_a_1[1] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[1] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I57_Y (.A(integral[8]), .B(
        \un1_next_int[8] ), .C(N345), .Y(N425));
    NOR3 inf_abs0_a_0_I_29 (.A(sr_new[7]), .B(sr_new[6]), .C(sr_new[8])
        , .Y(\DWACT_FINC_E_0[5] ));
    DFN1E0C0 \integ[23]  (.D(\un1_integ[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[23]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_2 (.A(
        ADD_26x26_fast_I206_un1_Y_0), .B(N522), .C(
        ADD_26x26_fast_I206_Y_1), .Y(ADD_26x26_fast_I206_Y_2));
    AO1 un1_integ_0_0_ADD_26x26_fast_I54_Y (.A(N344), .B(N348), .C(
        N347), .Y(N422));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I131_Y (.A(N405), .B(N401), .C(
        N462), .Y(N508));
    XNOR2 inf_abs0_a_0_I_26 (.A(sr_new[9]), .B(N_5), .Y(
        \inf_abs0_a_0[9] ));
    NOR3B inf_abs1_a_1_I_19 (.A(\DWACT_FINC_E[2] ), .B(
        \DWACT_FINC_E_0[0] ), .C(sr_old[6]), .Y(N_7));
    NOR3B inf_abs1_a_1_I_16 (.A(\DWACT_FINC_E[1] ), .B(
        \DWACT_FINC_E_0[0] ), .C(sr_old[5]), .Y(N_8));
    AX1D un1_integ_0_0_ADD_26x26_fast_I254_Y (.A(I205_un1_Y), .B(
        ADD_26x26_fast_I205_Y_3), .C(ADD_26x26_fast_I254_Y_0), .Y(
        \un1_integ[24] ));
    DFN1E0C0 \integ[19]  (.D(\un1_integ[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[19]));
    OR2 \state_RNIK2IJ2[1]  (.A(\un18_next_int_m[0] ), .B(
        \inf_abs1_m[0] ), .Y(\un1_next_int_iv_0[0] ));
    NOR2 inf_abs0_a_0_I_15 (.A(sr_new[3]), .B(sr_new[4]), .Y(
        \DWACT_FINC_E_0[1] ));
    MX2 \inf_abs1[8]  (.A(sr_old[8]), .B(\inf_abs1_a_1[8] ), .S(
        sr_old[12]), .Y(\inf_abs1[8]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I161_un1_Y (.A(N486), .B(N493), 
        .Y(I161_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I117_Y (.A(N439), .B(N435), .Y(
        N488));
    DFN1E0C0 \integ[17]  (.D(\un1_integ[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[17]));
    XOR2 inf_abs0_a_0_I_5 (.A(sr_new[0]), .B(sr_new[1]), .Y(
        \inf_abs0_a_0[1] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I33_Y (.A(integral[20]), .B(
        integral[21]), .C(\un1_next_int_0_iv_0[13] ), .Y(N401));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I255_Y_0 (.A(integral[25]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I255_Y_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I127_Y_0 (.A(integral[23]), .B(
        integral[22]), .C(\un1_next_int_0_iv[13] ), .Y(
        ADD_26x26_fast_I127_Y_0));
    OR3 \state_RNIN203C[0]  (.A(\inf_abs0_m[10] ), .B(
        \un1_next_int_iv_0[10] ), .C(\un2_next_int_m[10] ), .Y(
        \un1_next_int[10] ));
    DFN1E0C0 \integ[14]  (.D(\un1_integ[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[14]));
    XNOR2 inf_abs0_a_0_I_17 (.A(sr_new[6]), .B(N_8_0), .Y(
        \inf_abs0_a_0[6] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I87_Y (.A(N405), .B(N409), .Y(
        N458));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y_0 (.A(\integ[2]_net_1 ), 
        .B(\un1_next_int[2] ), .Y(ADD_26x26_fast_I232_Y_0));
    OR2 \state_RNI25NA4[0]  (.A(\un1_next_int_iv_1[0] ), .B(
        \un2_next_int_m[0] ), .Y(\un1_next_int[0] ));
    NOR2B \state_RNILBKG2[0]  (.A(\inf_abs0[6]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[6] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I84_Y (.A(N406), .B(I80_un1_Y), 
        .Y(N455));
    AO1 un1_integ_0_0_ADD_26x26_fast_I154_Y (.A(N485), .B(N478), .C(
        N477), .Y(N531));
    MX2 \inf_abs1[11]  (.A(sr_old[11]), .B(\inf_abs1_a_1[11] ), .S(
        sr_old[12]), .Y(\inf_abs1[11]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I11_G0N (.A(\un1_next_int[11] ), 
        .B(integral[11]), .Y(N350));
    NOR3B \state_RNI72R02[0]  (.A(sr_new_1_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[4]_net_1 ), .Y(\un2_next_int_m[4] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I140_Y (.A(N471), .B(N464), .C(
        N463), .Y(N517));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I149_Y (.A(N419), .B(N423), .C(
        N480), .Y(N526));
    NOR3B \state_RNISNFQ2[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[9] ), .Y(\un2_next_int_m[9] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I158_Y (.A(N489), .B(N482), .C(
        N481), .Y(N535));
    OR2 \state_RNIVTVR4[0]  (.A(\un1_next_int_iv_1[1] ), .B(
        \un2_next_int_m[1] ), .Y(\un1_next_int[1] ));
    OR2 \state_RNIRJ4F3[0]  (.A(\un1_next_int_iv_0[0] ), .B(
        \inf_abs0_m[0] ), .Y(\un1_next_int_iv_1[0] ));
    OR2 \state_RNIOMUD1_0[1]  (.A(next_int_1_sqmuxa), .B(
        next_int_0_sqmuxa_1), .Y(\un1_next_int_0_iv[13] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I249_Y_0 (.A(integral[19]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I249_Y_0));
    DFN1E0C0 \integ[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[25]));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I247_Y_0 (.A(integral[17]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I247_Y_0));
    XA1A \state_RNIJ18C5[1]  (.A(sr_old[12]), .B(\inf_abs1[8]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[8] ));
    OR3 \state_RNIAS3J4[1]  (.A(\inf_abs1_m[3] ), .B(
        \un18_next_int_m[3] ), .C(\inf_abs0_m[3] ), .Y(
        \un1_next_int_iv_1[3] ));
    MX2 \inf_abs1[6]  (.A(sr_old[6]), .B(\inf_abs1_a_1[6] ), .S(
        sr_old[12]), .Y(\inf_abs1[6]_net_1 ));
    NOR3 inf_abs0_a_0_I_33 (.A(sr_new[10]), .B(sr_new[9]), .C(
        sr_new[11]), .Y(\DWACT_FINC_E[7] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y_0 (.A(\integ[0]_net_1 ), 
        .B(N_3), .Y(ADD_26x26_fast_I230_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I64_un1_Y (.A(N329), .B(N333), 
        .Y(I64_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I242_Y (.A(N527), .B(I191_un1_Y), 
        .C(ADD_26x26_fast_I242_Y_0), .Y(\un1_integ[12] ));
    NOR3B \state_RNI5FMJ2[0]  (.A(sr_new_1_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[6]_net_1 ), .Y(\un2_next_int_m[6] ));
    XNOR2 inf_abs0_a_0_I_20 (.A(sr_new[7]), .B(N_7_0), .Y(
        \inf_abs0_a_0[7] ));
    NOR3B \state_RNI7HIR[0]  (.A(\state[0]_net_1 ), .B(sr_new_1_0), .C(
        sr_new[0]), .Y(\un2_next_int_m[0] ));
    DFN1E0C0 \integ[11]  (.D(\un1_integ[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[11]));
    MX2 \inf_abs0[8]  (.A(sr_new[8]), .B(\inf_abs0_a_0[8] ), .S(
        sr_new_1_0), .Y(\inf_abs0[8]_net_1 ));
    DFN1E0C0 \integ[16]  (.D(\un1_integ[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[16]));
    XNOR2 inf_abs1_a_1_I_28 (.A(sr_old[10]), .B(N_4), .Y(
        \inf_abs1_a_1[10] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I211_Y_1 (.A(
        ADD_26x26_fast_I211_un1_Y_0), .B(N531), .C(
        ADD_26x26_fast_I211_Y_1_0), .Y(ADD_26x26_fast_I211_Y_1));
    NOR3 inf_abs1_a_1_I_10 (.A(sr_old[1]), .B(sr_old[0]), .C(sr_old[2])
        , .Y(\DWACT_FINC_E_0[0] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I254_Y_0 (.A(integral[24]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I254_Y_0));
    OR2 \state_RNIVSL46[0]  (.A(\un1_next_int_iv_1[3] ), .B(
        \un2_next_int_m[3] ), .Y(\un1_next_int[3] ));
    MX2B un1_next_int_0_sqmuxa_0__m2 (.A(sr_new_1_0), .B(sr_old[12]), 
        .S(\state[1]_net_1 ), .Y(N_3));
    AO1 un1_integ_0_0_ADD_26x26_fast_I96_Y (.A(N418), .B(N415), .C(
        N414), .Y(N467));
    XA1A \state_RNI0R6I4[1]  (.A(sr_old[12]), .B(\inf_abs1[6]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[6] ));
    MX2 \inf_abs0[10]  (.A(sr_new[10]), .B(\inf_abs0_a_0[10] ), .S(
        sr_new_0_0), .Y(\inf_abs0[10]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I2_G0N (.A(\un1_next_int[2] ), 
        .B(\integ[2]_net_1 ), .Y(N323));
    AO1 un1_integ_0_0_ADD_26x26_fast_I114_Y (.A(N436), .B(N433), .C(
        N432), .Y(N485));
    OA1 un1_integ_0_0_ADD_26x26_fast_I189_un1_Y (.A(N485), .B(
        I161_un1_Y), .C(N524), .Y(I189_un1_Y));
    NOR2 inf_abs0_a_0_I_21 (.A(sr_new[6]), .B(sr_new[7]), .Y(
        \DWACT_FINC_E_0[3] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I147_Y (.A(N478), .B(N470), .Y(
        N524));
    DFN1E0C0 \integ[9]  (.D(\un1_integ[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(integral[9]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I242_Y_0 (.A(
        \un2_next_int_m[12] ), .B(\un1_next_int_iv_0[12] ), .C(
        integral[12]), .Y(ADD_26x26_fast_I242_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I235_Y (.A(N487), .B(I162_un1_Y), 
        .C(ADD_26x26_fast_I235_Y_0), .Y(\un1_integ[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I212_Y_0 (.A(N533), .B(N518), .C(
        N517), .Y(ADD_26x26_fast_I212_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I63_Y (.A(integral[6]), .B(
        \un1_next_int[6] ), .C(N333), .Y(N431));
    NOR2A inf_abs1_a_1_I_11 (.A(\DWACT_FINC_E_0[0] ), .B(sr_old[3]), 
        .Y(N_10_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I118_Y (.A(N440), .B(N437), .C(
        N436), .Y(N489));
    AX1D un1_integ_0_0_ADD_26x26_fast_I237_Y (.A(N483), .B(I160_un1_Y), 
        .C(ADD_26x26_fast_I237_Y_0), .Y(\un1_integ[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I133_Y (.A(N456), .B(N464), .Y(
        N510));
    NOR3B \state_RNINDFT2[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[10]_net_1 ), .Y(\un2_next_int_m[10] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I30_Y (.A(integral[22]), .B(
        integral[21]), .C(\un1_next_int_0_iv_0[13] ), .Y(N398));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I160_un1_Y (.A(N484), .B(N491), 
        .Y(I160_un1_Y));
    DFN1E0C0 \integ[22]  (.D(\un1_integ[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[22]));
    NOR3 inf_abs1_a_1_I_8 (.A(sr_old[1]), .B(sr_old[0]), .C(sr_old[2]), 
        .Y(N_11));
    AO1B un1_integ_0_0_ADD_26x26_fast_I43_Y (.A(integral[16]), .B(
        integral[15]), .C(\un1_next_int_0_iv_0[13] ), .Y(N411));
    NOR3C \state_RNIA1P91[1]  (.A(sr_old[0]), .B(\state[1]_net_1 ), .C(
        sr_old[12]), .Y(\inf_abs1_m[0] ));
    DFN1E0C0 \integ_0[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral_0_0));
    OR2 \state_RNIFPPM7[0]  (.A(\un1_next_int_iv_1[4] ), .B(
        \un2_next_int_m[4] ), .Y(\un1_next_int[4] ));
    DFN1E0C0 \integ[1]  (.D(\un1_integ[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(\integ[1]_net_1 ));
    OR2 \state_RNI8NUL5[1]  (.A(\un1_next_int_iv_0[4] ), .B(
        \inf_abs0_m[4] ), .Y(\un1_next_int_iv_1[4] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I35_Y (.A(integral[19]), .B(
        integral[20]), .C(\un1_next_int_0_iv_0[13] ), .Y(N403));
    NOR2B \state_RNI37QG2[1]  (.A(\inf_abs1_a_1[3] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[3] ));
    NOR2B inf_abs0_a_0_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I53_Y (.A(N348), .B(N351), .Y(
        N421));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I91_Y (.A(N409), .B(N413), .Y(
        N462));
    AX1D un1_integ_0_0_ADD_26x26_fast_I250_Y (.A(I178_un1_Y), .B(
        ADD_26x26_fast_I209_Y_1), .C(ADD_26x26_fast_I250_Y_0), .Y(
        \un1_integ[20] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I240_Y_0 (.A(integral[10]), .B(
        \un1_next_int[10] ), .Y(ADD_26x26_fast_I240_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I60_un1_Y (.A(N335), .B(N339), 
        .Y(I60_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_0 (.A(N467), .B(N460), .C(
        N459), .Y(ADD_26x26_fast_I210_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I71_Y (.A(\integ[2]_net_1 ), .B(
        \un1_next_int[2] ), .C(N321), .Y(N439));
    DFN1E0C0 \integ[20]  (.D(\un1_integ[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[20]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I244_Y (.A(N523), .B(I189_un1_Y), 
        .C(ADD_26x26_fast_I244_Y_0), .Y(\un1_integ[14] ));
    NOR3 inf_abs1_a_1_I_29 (.A(sr_old[7]), .B(sr_old[6]), .C(sr_old[8])
        , .Y(\DWACT_FINC_E[5] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I207_Y_1 (.A(N404), .B(N400), .C(
        N461), .Y(ADD_26x26_fast_I207_Y_1));
    OR2 un1_integ_0_0_ADD_26x26_fast_I106_Y (.A(I106_un1_Y), .B(N424), 
        .Y(N477));
    NOR2B \state_RNIUKGO[0]  (.A(sr_new[7]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[7] ));
    XNOR2 inf_abs0_a_0_I_32 (.A(sr_new[11]), .B(N_3_1), .Y(
        \inf_abs0_a_0[11] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_1 (.A(
        ADD_26x26_fast_I208_un1_Y_0), .B(N526), .C(
        ADD_26x26_fast_I208_Y_0), .Y(ADD_26x26_fast_I208_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I102_Y (.A(N424), .B(N421), .C(
        N420), .Y(N473));
    AX1D un1_integ_0_0_ADD_26x26_fast_I251_Y (.A(I176_un1_Y), .B(
        ADD_26x26_fast_I208_Y_1), .C(ADD_26x26_fast_I251_Y_0), .Y(
        \un1_integ[21] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I121_un1_Y (.A(N441), .B(
        \un1_next_int[0] ), .Y(I121_un1_Y));
    XNOR2 inf_abs1_a_1_I_26 (.A(sr_old[9]), .B(N_5_0), .Y(
        \inf_abs1_a_1[9] ));
    DFN1E0C0 \integ[18]  (.D(\un1_integ[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[18]));
    INV \integ_RNI07B1[24]  (.A(integral[24]), .Y(integral_i[24]));
    OR2 un1_integ_0_0_ADD_26x26_fast_I4_P0N (.A(\un1_next_int[4] ), .B(
        \integ[4]_net_1 ), .Y(N330));
    NOR3A \state_RNIF6P91[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .C(sr_old[5]), .Y(\un18_next_int_m[5] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I144_Y (.A(I144_un1_Y), .B(N467), 
        .Y(N521));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_0 (.A(N465), .B(N458), .C(
        N457), .Y(ADD_26x26_fast_I209_Y_0));
    OR3 \state_RNIQLHM9[0]  (.A(\inf_abs0_m[6] ), .B(
        \un1_next_int_iv_0[6] ), .C(\un2_next_int_m[6] ), .Y(
        \un1_next_int[6] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I148_Y (.A(I148_un1_Y), .B(N471), 
        .Y(N525));
    XA1A \state_RNIO6T66[1]  (.A(sr_old[12]), .B(\inf_abs1[10]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[10] ));
    XA1A \state_RNISQ7K6[1]  (.A(sr_old[12]), .B(\inf_abs1[11]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[11] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I60_Y (.A(I60_un1_Y), .B(N338), 
        .Y(N428));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y (.A(
        ADD_26x26_fast_I232_Y_0), .B(N493), .Y(\un1_integ[2] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I204_Y_2 (.A(N398), .B(
        ADD_26x26_fast_I204_Y_0), .C(N455), .Y(ADD_26x26_fast_I204_Y_2)
        );
    DFN1C0 \state[1]  (.D(\state_RNO_6[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[1]_net_1 ));
    XNOR2 inf_abs0_a_0_I_23 (.A(sr_new[8]), .B(N_6_0), .Y(
        \inf_abs0_a_0[8] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I110_un1_Y (.A(N432), .B(N429), 
        .Y(I110_un1_Y));
    NOR3A inf_abs1_a_1_I_13 (.A(\DWACT_FINC_E_0[0] ), .B(sr_old[3]), 
        .C(sr_old[4]), .Y(N_9));
    OA1 un1_integ_0_0_ADD_26x26_fast_I9_G0N (.A(\un2_next_int_m[9] ), 
        .B(\un1_next_int_iv_1[9] ), .C(integral[9]), .Y(N344));
    OA1B un1_integ_0_0_ADD_26x26_fast_I40_Y (.A(integral[17]), .B(
        integral[16]), .C(\un1_next_int_0_iv_0[13] ), .Y(N408));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I65_Y (.A(N333), .B(N330), .Y(
        N433));
    OA1 un1_integ_0_0_ADD_26x26_fast_I207_un1_Y_0 (.A(N485), .B(
        I161_un1_Y), .C(N508), .Y(ADD_26x26_fast_I207_un1_Y_0));
    NOR3 inf_abs0_a_0_I_8 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2]), 
        .Y(N_11_0));
    NOR3A \state_RNIC3P91[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .C(sr_old[2]), .Y(\un18_next_int_m[2] ));
    AND3 inf_abs1_a_1_I_30 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E_0[6] ));
    XNOR2 inf_abs0_a_0_I_35 (.A(sr_new[12]), .B(N_2), .Y(
        \inf_abs0_a_0[12] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I178_un1_Y (.A(N512), .B(N527), 
        .Y(I178_un1_Y));
    AO1B un1_integ_0_0_ADD_26x26_fast_I45_Y (.A(integral[15]), .B(
        integral[14]), .C(\un1_next_int_0_iv_0[13] ), .Y(N413));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I137_Y (.A(N419), .B(N415), .C(
        N460), .Y(N514));
    XNOR2 inf_abs0_a_0_I_9 (.A(sr_new[3]), .B(N_11_0), .Y(
        \inf_abs0_a_0[3] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I3_P0N (.A(\un1_next_int[3] ), .B(
        \integ[3]_net_1 ), .Y(N327));
    NOR2B \state_RNO[0]  (.A(N_46_1), .B(calc_int), .Y(
        \state_RNO_5[0] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I50_Y (.A(N350), .B(N354), .C(
        N353), .Y(N418));
    AO1 un1_integ_0_0_ADD_26x26_fast_I204_Y_3 (.A(N502), .B(N517), .C(
        ADD_26x26_fast_I204_Y_2), .Y(ADD_26x26_fast_I204_Y_3));
    XNOR2 inf_abs1_a_1_I_20 (.A(sr_old[7]), .B(N_7), .Y(
        \inf_abs1_a_1[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I74_un1_Y (.A(N318), .B(
        \un1_next_int[0] ), .Y(I74_un1_Y));
    XA1A \state_RNIHO5O3[1]  (.A(sr_old[12]), .B(\inf_abs1[4]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[4] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I36_Y (.A(integral[18]), .B(
        integral[19]), .C(\un1_next_int_0_iv_0[13] ), .Y(N404));
    NOR3A inf_abs1_a_1_I_31 (.A(\DWACT_FINC_E_0[6] ), .B(sr_old[9]), 
        .C(sr_old[10]), .Y(N_3_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I0_P0N (.A(N_3), .B(
        \integ[0]_net_1 ), .Y(N318));
    NOR2B \state_RNI0NGO[0]  (.A(sr_new[9]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[9] ));
    NOR2 inf_abs1_a_1_I_6 (.A(sr_old[0]), .B(sr_old[1]), .Y(N_12_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I55_Y (.A(N345), .B(N348), .Y(
        N423));
    OA1 un1_integ_0_0_ADD_26x26_fast_I205_un1_Y (.A(N535), .B(
        I195_un1_Y), .C(ADD_26x26_fast_I205_un1_Y_0), .Y(I205_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I163_un1_Y (.A(N490), .B(
        \un1_next_int[0] ), .Y(I163_un1_Y));
    OR3 \state_RNIHJQJC[0]  (.A(\inf_abs0_m[11] ), .B(
        \un1_next_int_iv_0[11] ), .C(\un2_next_int_m[11] ), .Y(
        \un1_next_int[11] ));
    NOR3A \state_RNIB2P91[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .C(sr_old[1]), .Y(\un18_next_int_m[1] ));
    NOR2 inf_abs1_a_1_I_21 (.A(sr_old[6]), .B(sr_old[7]), .Y(
        \DWACT_FINC_E[3] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I206_Y_1 (.A(N398), .B(I80_un1_Y), 
        .C(N459), .Y(ADD_26x26_fast_I206_Y_1));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I5_G0N (.A(\un1_next_int[5] ), 
        .B(\integ[5]_net_1 ), .Y(N332));
    NOR2B \state_RNIFPP32[1]  (.A(\inf_abs1_a_1[2] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[2] ));
    INV \integ_RNI18B1[25]  (.A(integral[25]), .Y(integral_i[25]));
    AND3 inf_abs0_a_0_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(
        \DWACT_FINC_E[4] ));
    DFN1E0C0 \integ[7]  (.D(\un1_integ[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(integral[7]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_2 (.A(
        ADD_26x26_fast_I207_un1_Y_0), .B(N524), .C(
        ADD_26x26_fast_I207_Y_1), .Y(ADD_26x26_fast_I207_Y_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I4_G0N (.A(\un1_next_int[4] ), 
        .B(\integ[4]_net_1 ), .Y(N329));
    NOR2B \state_RNIPFGO[0]  (.A(sr_new[2]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[2] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I206_un1_Y_0 (.A(N483), .B(
        I160_un1_Y), .C(N506), .Y(ADD_26x26_fast_I206_un1_Y_0));
    XNOR2 inf_abs1_a_1_I_14 (.A(sr_old[5]), .B(N_9), .Y(
        \inf_abs1_a_1[5] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I234_Y (.A(N489), .B(I163_un1_Y), 
        .C(ADD_26x26_fast_I234_Y_0), .Y(\un1_integ[4] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I205_Y_2 (.A(N400), .B(
        ADD_26x26_fast_I205_Y_0), .C(N457), .Y(ADD_26x26_fast_I205_Y_2)
        );
    NOR2B un1_integ_0_0_ADD_26x26_fast_I174_un1_Y (.A(N508), .B(N523), 
        .Y(I174_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I162_un1_Y (.A(N488), .B(N442), 
        .Y(I162_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I240_Y (.A(N531), .B(I193_un1_Y), 
        .C(ADD_26x26_fast_I240_Y_0), .Y(\un1_integ[10] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I156_Y (.A(N487), .B(N480), .C(
        N479), .Y(N533));
    OR2 \state_RNIOMUD1[1]  (.A(next_int_1_sqmuxa), .B(
        next_int_0_sqmuxa_1), .Y(\un1_next_int_0_iv_0[13] ));
    DFN1E0C0 \integ[8]  (.D(\un1_integ[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(integral[8]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I85_Y (.A(N407), .B(N403), .Y(
        N456));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I251_Y_0 (.A(integral[21]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I251_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I152_Y (.A(N483), .B(N476), .C(
        N475), .Y(N529));
    AND3 inf_abs0_a_0_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(N_6_0));
    OR3 un1_integ_0_0_ADD_26x26_fast_I9_P0N (.A(\un2_next_int_m[9] ), 
        .B(\un1_next_int_iv_1[9] ), .C(integral[9]), .Y(N345));
    OA1 un1_integ_0_0_ADD_26x26_fast_I208_un1_Y_0 (.A(N487), .B(
        I162_un1_Y), .C(N510), .Y(ADD_26x26_fast_I208_un1_Y_0));
    OR2 \state_RNIVT2P3[0]  (.A(\un1_next_int_iv_0[1] ), .B(
        \inf_abs0_m[1] ), .Y(\un1_next_int_iv_1[1] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I31_Y (.A(integral[21]), .B(
        integral[22]), .C(\un1_next_int_0_iv_0[13] ), .Y(N399));
    XNOR2 inf_abs1_a_1_I_12 (.A(sr_old[4]), .B(N_10_0), .Y(
        \inf_abs1_a_1[4] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I235_Y_0 (.A(\integ[5]_net_1 ), 
        .B(\un1_next_int[5] ), .Y(ADD_26x26_fast_I235_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I56_un1_Y (.A(integral[8]), .B(
        \un1_next_int[8] ), .C(N345), .Y(I56_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I241_Y (.A(N529), .B(I192_un1_Y), 
        .C(ADD_26x26_fast_I241_Y_0), .Y(\un1_integ[11] ));
    NOR3A \state_RNIJAP91[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .C(sr_old[9]), .Y(\un18_next_int_m[9] ));
    NOR3 inf_abs0_a_0_I_18 (.A(sr_new[4]), .B(sr_new[3]), .C(sr_new[5])
        , .Y(\DWACT_FINC_E_0[2] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I11_P0N (.A(\un1_next_int[11] ), 
        .B(integral[11]), .Y(N351));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I243_Y_0 (.A(integral[13]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I243_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I105_Y (.A(N427), .B(N423), .Y(
        N476));
    AO1 un1_integ_0_0_ADD_26x26_fast_I213_Y_0 (.A(N535), .B(N520), .C(
        N519), .Y(ADD_26x26_fast_I213_Y_0));
    MX2 \inf_abs0[11]  (.A(sr_new[11]), .B(\inf_abs0_a_0[11] ), .S(
        sr_new_0_0), .Y(\inf_abs0[11]_net_1 ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I238_Y_0 (.A(integral[8]), .B(
        \un1_next_int[8] ), .Y(ADD_26x26_fast_I238_Y_0));
    NOR3A \state_RNIA1P91_0[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .C(sr_old[0]), .Y(\un18_next_int_m[0] ));
    XOR2 inf_abs1_a_1_I_5 (.A(sr_old[0]), .B(sr_old[1]), .Y(
        \inf_abs1_a_1[1] ));
    NOR3B \state_RNIE5702[0]  (.A(sr_new_1_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[5] ), .Y(\un2_next_int_m[5] ));
    NOR3A \state_RNID4P91[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .C(sr_old[3]), .Y(\un18_next_int_m[3] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I66_Y (.A(N326), .B(N330), .C(
        N329), .Y(N434));
    AX1D un1_integ_0_0_ADD_26x26_fast_I248_Y (.A(
        ADD_26x26_fast_I211_Y_1), .B(ADD_26x26_fast_I211_Y_0), .C(
        ADD_26x26_fast_I248_Y_0), .Y(\un1_integ[18] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I99_Y (.A(N417), .B(N421), .Y(
        N470));
    OR2 un1_integ_0_0_ADD_26x26_fast_I92_Y (.A(N414), .B(N410), .Y(
        N463));
    OA1 un1_integ_0_0_ADD_26x26_fast_I191_un1_Y (.A(N489), .B(
        I163_un1_Y), .C(N528), .Y(I191_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I72_Y (.A(N317), .B(N321), .C(
        N320), .Y(N440));
    OR3 \state_RNI3G717[1]  (.A(\inf_abs0_m[9] ), .B(
        \un18_next_int_m[9] ), .C(\inf_abs1_m[9] ), .Y(
        \un1_next_int_iv_1[9] ));
    NOR2B \state_RNIGETU4[1]  (.A(\inf_abs1_a_1[9] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[9] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I46_Y (.A(integral[13]), .B(
        integral[14]), .C(\un1_next_int_0_iv_0[13] ), .Y(N414));
    NOR2 \state_RNI94SU[0]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 )
        , .Y(N_46_1));
    NOR3 inf_abs1_a_1_I_33 (.A(sr_old[10]), .B(sr_old[9]), .C(
        sr_old[11]), .Y(\DWACT_FINC_E_0[7] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I116_Y (.A(N438), .B(N435), .C(
        N434), .Y(N487));
    OR2 \state_RNI7FI03[1]  (.A(\un18_next_int_m[1] ), .B(
        \inf_abs1_m[1] ), .Y(\un1_next_int_iv_0[1] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I112_Y (.A(N434), .B(N431), .C(
        N430), .Y(N483));
    NOR2A inf_abs0_a_0_I_25 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .Y(
        N_5));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I213_un1_Y_0 (.A(N482), .B(N490)
        , .C(\un1_next_int[0] ), .Y(ADD_26x26_fast_I213_un1_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I210_un1_Y (.A(N514), .B(N491), 
        .C(N530), .Y(I210_un1_Y));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y_0 (.A(\integ[4]_net_1 ), 
        .B(\un1_next_int[4] ), .Y(ADD_26x26_fast_I234_Y_0));
    NOR3A inf_abs0_a_0_I_27 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .C(
        sr_new[9]), .Y(N_4_0));
    
endmodule


module error_calc_13s_12s_4_2(
       cur_error,
       LED_5_i_0,
       LED_5,
       average,
       calc_error,
       n_rst_c,
       clk_c
    );
output [12:0] cur_error;
input  LED_5_i_0;
input  [7:0] LED_5;
input  [6:2] average;
input  calc_error;
input  n_rst_c;
input  clk_c;

    wire N_40, N_38, GND, VCC;
    
    AX1B un2_diffreg_1_m37 (.A(LED_5[5]), .B(LED_5[6]), .C(LED_5[7]), 
        .Y(N_38));
    DFN1E1C0 \diffreg[3]  (.D(average[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[3]));
    XNOR2 un2_diffreg_1_m39 (.A(LED_5[6]), .B(LED_5[5]), .Y(N_40));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \diffreg[7]  (.D(LED_5[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[7]));
    DFN1E1C0 \diffreg[1]  (.D(average[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[1]));
    DFN1E1C0 \diffreg[12]  (.D(N_38), .CLK(clk_c), .CLR(n_rst_c), .E(
        calc_error), .Q(cur_error[12]));
    DFN1E1C0 \diffreg[11]  (.D(N_40), .CLK(clk_c), .CLR(n_rst_c), .E(
        calc_error), .Q(cur_error[11]));
    GND GND_i (.Y(GND));
    DFN1E1C0 \diffreg[9]  (.D(LED_5[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[9]));
    DFN1E1C0 \diffreg[8]  (.D(LED_5[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[8]));
    DFN1E1C0 \diffreg[6]  (.D(LED_5[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[6]));
    DFN1E1C0 \diffreg[10]  (.D(LED_5_i_0), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[10]));
    DFN1E1C0 \diffreg[5]  (.D(LED_5[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[5]));
    DFN1E1C0 \diffreg[4]  (.D(average[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[4]));
    DFN1E1C0 \diffreg[2]  (.D(average[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[2]));
    DFN1E1C0 \diffreg[0]  (.D(average[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[0]));
    
endmodule


module derivative_calc_13s_4_2(
       derivative_0,
       sr_prev,
       sr_new,
       sr_new_0_0,
       deriv_enable,
       n_rst_c,
       clk_c
    );
output derivative_0;
input  [12:0] sr_prev;
input  [11:0] sr_new;
input  sr_new_0_0;
input  deriv_enable;
input  n_rst_c;
input  clk_c;

    wire SUB_13x13_medium_area_I49_Y_1, N208, N176, 
        SUB_13x13_medium_area_I49_Y_0, 
        SUB_13x13_medium_area_I26_un1_Y_0, 
        SUB_13x13_medium_area_I49_un1_Y_1, 
        SUB_13x13_medium_area_I49_un1_Y_0, N_15, 
        SUB_13x13_medium_area_I42_Y_1, N218, N180, 
        SUB_13x13_medium_area_I42_Y_0, 
        SUB_13x13_medium_area_I30_un1_Y_0, 
        SUB_13x13_medium_area_I42_un1_Y_1, N_9, N_7, 
        SUB_13x13_medium_area_I41_Y_0, 
        SUB_13x13_medium_area_I34_un1_Y_0, 
        SUB_13x13_medium_area_I41_un1_Y_0, N_5, 
        SUB_13x13_medium_area_I28_un1_Y_0, 
        SUB_13x13_medium_area_I32_un1_Y_0, N212, N222, N_24, N226, 
        N204, N185, N_21, N_13, GND, VCC;
    
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I34_un1_Y_0 (.A(
        sr_new[1]), .B(sr_prev[1]), .Y(
        SUB_13x13_medium_area_I34_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y_0 (.A(
        SUB_13x13_medium_area_I30_un1_Y_0), .B(sr_new[6]), .C(
        sr_prev[6]), .Y(SUB_13x13_medium_area_I42_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I15_S (.A(sr_prev[2]), 
        .B(sr_new[2]), .Y(N_5));
    OR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I36_Y (.A(sr_prev[0]), 
        .B(sr_new[0]), .Y(N185));
    XNOR3 un2_deriv_out_0_0_SUB_13x13_medium_area_I82_Y (.A(sr_new_0_0)
        , .B(sr_prev[12]), .C(N226), .Y(N_24));
    VCC VCC_i (.Y(VCC));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I64_Y (.A(N204), .B(
        sr_new[11]), .C(sr_prev[11]), .Y(N226));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I41_Y_0 (.A(
        SUB_13x13_medium_area_I34_un1_Y_0), .B(sr_new[2]), .C(
        sr_prev[2]), .Y(SUB_13x13_medium_area_I41_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I19_S (.A(sr_prev[6]), 
        .B(sr_new[6]), .Y(N_13));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I28_Y (.A(
        SUB_13x13_medium_area_I28_un1_Y_0), .B(sr_new[8]), .C(
        sr_prev[8]), .Y(N208));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y_1 (.A(N218), .B(
        N180), .C(SUB_13x13_medium_area_I42_Y_0), .Y(
        SUB_13x13_medium_area_I42_Y_1));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I28_un1_Y_0 (.A(
        sr_new[7]), .B(sr_prev[7]), .Y(
        SUB_13x13_medium_area_I28_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y_0 (.A(
        SUB_13x13_medium_area_I26_un1_Y_0), .B(sr_new[10]), .C(
        sr_prev[10]), .Y(SUB_13x13_medium_area_I49_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I20_S (.A(sr_prev[7]), 
        .B(sr_new[7]), .Y(N_15));
    DFN1E1C0 \deriv_out[12]  (.D(N_24), .CLK(clk_c), .CLR(n_rst_c), .E(
        deriv_enable), .Q(derivative_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I17_S (.A(sr_prev[4]), 
        .B(sr_new[4]), .Y(N_9));
    GND GND_i (.Y(GND));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I23_S (.A(sr_prev[10])
        , .B(sr_new[10]), .Y(N_21));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I26_un1_Y_0 (.A(
        sr_new[9]), .B(sr_prev[9]), .Y(
        SUB_13x13_medium_area_I26_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I32_Y (.A(
        SUB_13x13_medium_area_I32_un1_Y_0), .B(sr_new[4]), .C(
        sr_prev[4]), .Y(N218));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I30_un1_Y_0 (.A(
        sr_new[5]), .B(sr_prev[5]), .Y(
        SUB_13x13_medium_area_I30_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y (.A(
        SUB_13x13_medium_area_I49_un1_Y_1), .B(N212), .C(
        SUB_13x13_medium_area_I49_Y_1), .Y(N204));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I32_un1_Y_0 (.A(
        sr_new[3]), .B(sr_prev[3]), .Y(
        SUB_13x13_medium_area_I32_un1_Y_0));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I31_Y (.A(sr_new[5]), 
        .B(sr_prev[5]), .C(N_13), .Y(N180));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I41_un1_Y_0 (.A(
        sr_new[1]), .B(sr_prev[1]), .C(N_5), .Y(
        SUB_13x13_medium_area_I41_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y_1 (.A(N208), .B(
        N176), .C(SUB_13x13_medium_area_I49_Y_0), .Y(
        SUB_13x13_medium_area_I49_Y_1));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I16_S (.A(sr_prev[3]), 
        .B(sr_new[3]), .Y(N_7));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y (.A(
        SUB_13x13_medium_area_I42_un1_Y_1), .B(N222), .C(
        SUB_13x13_medium_area_I42_Y_1), .Y(N212));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I27_Y (.A(sr_new[9]), 
        .B(sr_prev[9]), .C(N_21), .Y(N176));
    NOR2B un2_deriv_out_0_0_SUB_13x13_medium_area_I49_un1_Y_1 (.A(
        SUB_13x13_medium_area_I49_un1_Y_0), .B(N176), .Y(
        SUB_13x13_medium_area_I49_un1_Y_1));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I49_un1_Y_0 (.A(
        sr_new[8]), .B(sr_prev[8]), .C(N_15), .Y(
        SUB_13x13_medium_area_I49_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I41_Y (.A(
        SUB_13x13_medium_area_I41_un1_Y_0), .B(N185), .C(
        SUB_13x13_medium_area_I41_Y_0), .Y(N222));
    NOR3A un2_deriv_out_0_0_SUB_13x13_medium_area_I42_un1_Y_1 (.A(N180)
        , .B(N_9), .C(N_7), .Y(SUB_13x13_medium_area_I42_un1_Y_1));
    
endmodule


module pwm_tx_400s_32s_13s_10_222s_45s(
       off_div,
       act_ctl_5_i,
       act_ctl_5_1,
       act_ctl_5_0,
       pwm_chg_0,
       pwm_chg,
       n_rst_c,
       clk_c,
       act_ctl_5_7,
       act_ctl_5_6,
       act_ctl_5_8,
       act_ctl_5_4,
       primary_5_c
    );
input  [31:0] off_div;
input  act_ctl_5_i;
input  act_ctl_5_1;
input  act_ctl_5_0;
input  pwm_chg_0;
input  pwm_chg;
input  n_rst_c;
input  clk_c;
input  act_ctl_5_7;
input  act_ctl_5_6;
input  act_ctl_5_8;
input  act_ctl_5_4;
output primary_5_c;

    wire N_400_0, I_140_6, I_140_5, \DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] , \DWACT_COMP0_E[1] , N_18, 
        I_20_6, \counter[7]_net_1 , N_20, I_23_9, \counter[8]_net_1 , 
        N_11, N_6, N_8, \DWACT_FDEC_E[0] , N_3, \DWACT_FDEC_E[2] , 
        N_16, N_14, \counter[6]_net_1 , N_2, \counter[2]_net_1 , 
        counter_m6_0_a2_7, counter_m6_0_a2_2, counter_m6_0_a2_1, 
        counter_m6_0_a2_6, \counter[16]_net_1 , \counter[18]_net_1 , 
        counter_m6_0_a2_4, \counter[15]_net_1 , \counter[10]_net_1 , 
        \counter[17]_net_1 , \counter[13]_net_1 , \counter[14]_net_1 , 
        \counter[11]_net_1 , \counter[12]_net_1 , counter_c18, 
        \counter[9]_net_1 , counter_c8, counter_n31, 
        \counter[31]_net_1 , counter_63_0, cur_pwm_RNIQQ9OA2_0_net_1, 
        \counter[30]_net_1 , counter_c29, counter_n30, counter_n29, 
        \counter[29]_net_1 , counter_c28, counter_n28, counter_n28_tz, 
        \counter[27]_net_1 , counter_c26, \counter[28]_net_1 , 
        counter_n27, counter_n26, counter_n26_tz, \counter[25]_net_1 , 
        counter_c24, \counter[26]_net_1 , counter_n25, counter_n24, 
        counter_n24_tz, \counter[23]_net_1 , counter_c22, 
        \counter[24]_net_1 , counter_n23, counter_n22, counter_n22_tz, 
        \counter[21]_net_1 , counter_c20, \counter[22]_net_1 , 
        counter_n21, counter_n20, counter_n20_tz, \counter[19]_net_1 , 
        \counter[20]_net_1 , counter_n19, counter_n18, counter_c17, 
        counter_n17, counter_c16, counter_n16, counter_c15, 
        counter_n15, counter_c14, counter_n14, counter_c13, 
        counter_n13, counter_c12, counter_n12, counter_c11, 
        counter_n11, counter_c10, counter_n10, counter_n10_tz, 
        counter_n9, counter_n8, counter_n8_tz, counter_c6, counter_n7, 
        counter_n6, counter_n6_tz, \counter[5]_net_1 , counter_c4, 
        counter_n5, counter_n4, counter_n4_tz, \counter[3]_net_1 , 
        counter_c2, \counter[4]_net_1 , counter_n3, counter_n2, 
        counter_n2_tz, \counter[1]_net_1 , \counter[0]_net_1 , 
        \off_time[0] , \off_reg[0]_net_1 , \off_time[1] , 
        \off_reg[1]_net_1 , \off_time[2] , \off_reg[2]_net_1 , 
        \off_time[3] , \off_reg[3]_net_1 , \off_time[4] , 
        \off_reg[4]_net_1 , \off_time[6] , \off_reg[6]_net_1 , 
        \off_time[9] , \off_reg[9]_net_1 , \off_time[11] , 
        \off_reg[11]_net_1 , \off_time[13] , \off_reg[13]_net_1 , 
        \off_time[17] , \off_reg[17]_net_1 , \off_time[18] , 
        \off_reg[18]_net_1 , \off_time[20] , \off_reg[20]_net_1 , 
        \off_time[21] , \off_reg[21]_net_1 , \off_time[22] , 
        \off_reg[22]_net_1 , \off_time[25] , \off_reg[25]_net_1 , 
        \off_time[30] , \off_reg[30]_net_1 , \off_time[31] , 
        \off_reg[31]_net_1 , \off_time[14] , \off_reg[14]_net_1 , 
        \off_time[16] , \off_reg[16]_net_1 , \off_time[7] , 
        \off_reg[7]_net_1 , \off_time[5] , \off_reg[5]_net_1 , 
        \off_time[28] , \off_reg[28]_net_1 , \off_time[15] , 
        \off_reg[15]_net_1 , \off_time[26] , \off_reg[26]_net_1 , 
        \off_time[29] , \off_reg[29]_net_1 , \off_time[27] , 
        \off_reg[27]_net_1 , \off_time[24] , \off_reg[24]_net_1 , 
        \off_time[23] , \off_reg[23]_net_1 , \off_time[8] , 
        \off_reg[8]_net_1 , \off_time[12] , \off_reg[12]_net_1 , 
        \off_time[19] , \off_reg[19]_net_1 , \off_time[10] , 
        \off_reg[10]_net_1 , counter_n1, \counter_RNO_2[0] , 
        cur_pwm_RNO_2, \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] , N_4, N_21, N_17, N_13, 
        I_14_6, \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] , \DWACT_BL_EQUAL_0_E[3] , 
        \DWACT_BL_EQUAL_0_E[2] , \DWACT_BL_EQUAL_0_E[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] , \DWACT_COMP0_E_0[1] , 
        \DWACT_COMP0_E_0[2] , \DWACT_COMP0_E[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] , N_11_0, N_10, N_9, N_6_0, 
        N_8_0, N_7, N_5, N_2_0, N_3_0, N_4_0, N_21_0, N_20_0, N_19, 
        N_16_0, N_18_0, N_17_0, N_15, N_12, N_13_0, N_14_0, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] , 
        \DWACT_BL_EQUAL_0_E[4] , \DWACT_BL_EQUAL_0_E_0[3] , 
        \DWACT_BL_EQUAL_0_E_0[0] , \DWACT_BL_EQUAL_0_E[1] , 
        \DWACT_BL_EQUAL_0_E_0[2] , \DWACT_CMPLE_PO0_DWACT_COMP0_E[1] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[0] , N_31, N_30, N_29, N_26, 
        N_28, N_27, N_25, N_22, N_23, N_24, \ACT_LT4_E[3] , 
        \ACT_LT4_E[6] , \ACT_LT4_E[10] , \ACT_LT4_E[7] , 
        \ACT_LT4_E[8] , \ACT_LT4_E[5] , \ACT_LT4_E[4] , \ACT_LT4_E[0] , 
        \ACT_LT4_E[1] , \ACT_LT4_E[2] , \DWACT_BL_EQUAL_0_E_1[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] , 
        \DWACT_BL_EQUAL_0_E_1[0] , \DWACT_BL_EQUAL_0_E_0[1] , 
        \DWACT_BL_EQUAL_0_E_1[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] , 
        \DWACT_BL_EQUAL_0_E_2[0] , \DWACT_BL_EQUAL_0_E_1[1] , 
        \DWACT_BL_EQUAL_0_E_2[2] , \DWACT_BL_EQUAL_0_E_2[3] , 
        \DWACT_BL_EQUAL_0_E_0[4] , \DWACT_BL_EQUAL_0_E[5] , 
        \DWACT_BL_EQUAL_0_E[6] , \DWACT_BL_EQUAL_0_E[7] , 
        \DWACT_BL_EQUAL_0_E[8] , \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] , N_41, N_40, N_39, N_36, 
        N_38, N_37, N_35, N_32, N_33, N_34, \ACT_LT3_E[3] , 
        \ACT_LT3_E[4] , \ACT_LT3_E[5] , \ACT_LT3_E[0] , \ACT_LT3_E[1] , 
        \ACT_LT3_E[2] , \DWACT_BL_EQUAL_0_E_3[2] , 
        \DWACT_BL_EQUAL_0_E_2[1] , \DWACT_BL_EQUAL_0_E_3[0] , N_51, 
        N_50, N_49, N_46, N_48, N_47, N_45, N_42, N_43, N_44, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] , 
        \DWACT_BL_EQUAL_0_E_1[4] , \DWACT_BL_EQUAL_0_E_3[3] , 
        \DWACT_BL_EQUAL_0_E_4[0] , \DWACT_BL_EQUAL_0_E_3[1] , 
        \DWACT_BL_EQUAL_0_E_4[2] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] , 
        \DWACT_BL_EQUAL_0_E[12] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] , 
        \DWACT_BL_EQUAL_0_E_5[0] , \DWACT_BL_EQUAL_0_E_4[1] , 
        \DWACT_BL_EQUAL_0_E_5[2] , \DWACT_BL_EQUAL_0_E_4[3] , 
        \DWACT_BL_EQUAL_0_E_2[4] , \DWACT_BL_EQUAL_0_E_0[5] , 
        \DWACT_BL_EQUAL_0_E_0[6] , \DWACT_BL_EQUAL_0_E_0[7] , 
        \DWACT_BL_EQUAL_0_E_0[8] , \DWACT_BL_EQUAL_0_E[9] , 
        \DWACT_BL_EQUAL_0_E[10] , \DWACT_BL_EQUAL_0_E[11] , N_2_1, 
        N_5_0, GND, VCC;
    
    OR2 \off_reg_RNIR0RG[7]  (.A(\off_reg[7]_net_1 ), .B(act_ctl_5_8), 
        .Y(\off_time[7] ));
    DFN1C0 \counter[19]  (.D(counter_n19), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[19]_net_1 ));
    AND3 un1_counter_0_I_78 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] ));
    NOR3 un1_counter_2_0_I_17 (.A(\counter[20]_net_1 ), .B(
        \counter[19]_net_1 ), .C(\counter[21]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] ));
    XOR2 un1_act_ctl_I_23 (.A(act_ctl_5_4), .B(N_2_1), .Y(I_23_9));
    AND2A un1_counter_0_I_51 (.A(\off_time[26] ), .B(
        \counter[26]_net_1 ), .Y(\ACT_LT3_E[5] ));
    OR2 \off_reg_RNIQVQG[6]  (.A(\off_reg[6]_net_1 ), .B(act_ctl_5_8), 
        .Y(\off_time[6] ));
    DFN1E1C0 \off_reg[28]  (.D(off_div[28]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[28]_net_1 ));
    AX1C \counter_RNO_0[2]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .C(\counter[2]_net_1 ), .Y(counter_n2_tz));
    MX2C cur_pwm_RNIQQ9OA2_0 (.A(I_140_6), .B(I_140_5), .S(primary_5_c)
        , .Y(cur_pwm_RNIQQ9OA2_0_net_1));
    DFN1C0 \counter[28]  (.D(counter_n28), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[28]_net_1 ));
    XNOR2 un1_counter_0_I_73 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .Y(\DWACT_BL_EQUAL_0_E_2[2] ));
    OA1A un1_counter_0_I_136 (.A(N_6_0), .B(N_8_0), .C(N_7), .Y(N_11_0)
        );
    OA1A un1_counter_0_I_132 (.A(\counter[3]_net_1 ), .B(\off_time[3] )
        , .C(N_3_0), .Y(N_7));
    NOR2A \off_reg_RNI4NSC[11]  (.A(\off_reg[11]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[11] ));
    DFN1E1C0 \off_reg[15]  (.D(off_div[15]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[15]_net_1 ));
    DFN1E1C0 \off_reg[26]  (.D(off_div[26]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[26]_net_1 ));
    NOR3C \counter_RNI67V43[9]  (.A(\counter[9]_net_1 ), .B(counter_c8)
        , .C(counter_m6_0_a2_7), .Y(counter_c18));
    AND3 un1_counter_0_I_14 (.A(\DWACT_BL_EQUAL_0_E[9] ), .B(
        \DWACT_BL_EQUAL_0_E[10] ), .C(\DWACT_BL_EQUAL_0_E[11] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] ));
    XA1B \counter_RNO[11]  (.A(\counter[11]_net_1 ), .B(counter_c10), 
        .C(N_400_0), .Y(counter_n11));
    NOR3C \counter_RNISP2A4[24]  (.A(\counter[23]_net_1 ), .B(
        counter_c22), .C(\counter[24]_net_1 ), .Y(counter_c24));
    DFN1C0 \counter[29]  (.D(counter_n29), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[29]_net_1 ));
    DFN1E1C0 \off_reg[5]  (.D(off_div[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[5]_net_1 ));
    NOR3 un1_counter_2_0_I_77 (.A(\counter[12]_net_1 ), .B(
        \counter[10]_net_1 ), .C(\counter[11]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] ));
    XNOR2 un1_counter_0_I_82 (.A(\counter[15]_net_1 ), .B(
        \off_time[15] ), .Y(\DWACT_BL_EQUAL_0_E_1[0] ));
    DFN1C0 \counter[11]  (.D(counter_n11), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[11]_net_1 ));
    XNOR2 un1_counter_0_I_109 (.A(\counter[6]_net_1 ), .B(
        \off_time[6] ), .Y(\DWACT_BL_EQUAL_0_E[1] ));
    NOR2A \off_reg_RNICVSC[19]  (.A(\off_reg[19]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[19] ));
    NOR2A un1_counter_2_0_I_118 (.A(I_14_6), .B(\counter[5]_net_1 ), 
        .Y(N_14));
    OR2A un1_counter_0_I_103 (.A(\counter[14]_net_1 ), .B(
        \off_time[14] ), .Y(N_29));
    NOR2A \counter_RNO[28]  (.A(counter_n28_tz), .B(
        cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n28));
    XA1B \counter_RNO[15]  (.A(\counter[15]_net_1 ), .B(counter_c14), 
        .C(N_400_0), .Y(counter_n15));
    NOR3C \counter_RNIJ5FM4[26]  (.A(\counter[25]_net_1 ), .B(
        counter_c24), .C(\counter[26]_net_1 ), .Y(counter_c26));
    XNOR2 un1_counter_0_I_25 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .Y(\DWACT_BL_EQUAL_0_E_3[3] ));
    AND2 un1_counter_0_I_114 (.A(\DWACT_BL_EQUAL_0_E[4] ), .B(
        \DWACT_BL_EQUAL_0_E_0[3] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] ));
    XNOR2 un1_counter_0_I_11 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .Y(\DWACT_BL_EQUAL_0_E_4[3] ));
    NOR2B \counter_RNIDV9C[11]  (.A(\counter[11]_net_1 ), .B(
        \counter[12]_net_1 ), .Y(counter_m6_0_a2_1));
    OR3A un1_act_ctl_I_22 (.A(act_ctl_5_1), .B(\DWACT_FDEC_E[2] ), .C(
        \DWACT_FDEC_E[0] ), .Y(N_2_1));
    NOR2B \counter_RNI7G002[12]  (.A(counter_c11), .B(
        \counter[12]_net_1 ), .Y(counter_c12));
    OR2 \off_reg_RNIOTQG[4]  (.A(\off_reg[4]_net_1 ), .B(act_ctl_5_8), 
        .Y(\off_time[4] ));
    AX1C \counter_RNO_0[22]  (.A(\counter[21]_net_1 ), .B(counter_c20), 
        .C(\counter[22]_net_1 ), .Y(counter_n22_tz));
    XA1B \counter_RNO[7]  (.A(\counter[7]_net_1 ), .B(counter_c6), .C(
        N_400_0), .Y(counter_n7));
    OA1A un1_counter_2_0_I_125 (.A(N_16), .B(N_18), .C(N_17), .Y(N_21));
    DFN1E1C0 \off_reg[2]  (.D(off_div[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[2]_net_1 ));
    XNOR2 un1_counter_0_I_72 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .Y(\DWACT_BL_EQUAL_0_E_2[3] ));
    OA1 un1_counter_0_I_126 (.A(N_21_0), .B(N_20_0), .C(N_19), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] ));
    DFN1C0 \counter[6]  (.D(counter_n6), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[6]_net_1 ));
    AO1C un1_counter_0_I_122 (.A(\counter[7]_net_1 ), .B(\off_time[7] )
        , .C(N_12), .Y(N_18_0));
    XA1B \counter_RNO[31]  (.A(\counter[31]_net_1 ), .B(counter_63_0), 
        .C(cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n31));
    DFN1C0 \counter[21]  (.D(counter_n21), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[21]_net_1 ));
    AND2 un1_counter_0_I_20 (.A(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] ), .B(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] ), .Y(
        \DWACT_COMP0_E_0[1] ));
    OR2 un1_act_ctl_I_10 (.A(act_ctl_5_4), .B(act_ctl_5_4), .Y(
        \DWACT_FDEC_E[0] ));
    NOR2A \off_reg_RNI9SSC[16]  (.A(\off_reg[16]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[16] ));
    NOR2B \counter_RNI2NFI2[15]  (.A(counter_c14), .B(
        \counter[15]_net_1 ), .Y(counter_c15));
    DFN1C0 \counter[3]  (.D(counter_n3), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[3]_net_1 ));
    DFN1C0 \counter[2]  (.D(counter_n2), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[2]_net_1 ));
    AND3 un1_counter_0_I_45 (.A(\DWACT_BL_EQUAL_0_E_3[2] ), .B(
        \DWACT_BL_EQUAL_0_E_2[1] ), .C(\DWACT_BL_EQUAL_0_E_3[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] ));
    NOR2A \off_reg_RNI7U1E[31]  (.A(\off_reg[31]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[31] ));
    DFN1E1C0 \off_reg[23]  (.D(off_div[23]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[23]_net_1 ));
    NOR2A \counter_RNO[8]  (.A(counter_n8_tz), .B(
        cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n8));
    OA1A un1_counter_2_0_I_121 (.A(\counter[8]_net_1 ), .B(I_23_9), .C(
        N_13), .Y(N_17));
    XA1B \counter_RNO[13]  (.A(\counter[13]_net_1 ), .B(counter_c12), 
        .C(N_400_0), .Y(counter_n13));
    AO1C un1_counter_0_I_57 (.A(\off_time[20] ), .B(
        \counter[20]_net_1 ), .C(N_34), .Y(N_36));
    DFN1E1C0 \off_reg[9]  (.D(off_div[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[9]_net_1 ));
    XNOR2 un1_counter_0_I_26 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(\DWACT_BL_EQUAL_0_E_4[2] ));
    AX1C \counter_RNO_0[4]  (.A(\counter[3]_net_1 ), .B(counter_c2), 
        .C(\counter[4]_net_1 ), .Y(counter_n4_tz));
    AO1C un1_counter_0_I_35 (.A(\off_time[28] ), .B(
        \counter[28]_net_1 ), .C(N_44), .Y(N_46));
    AO1 un1_counter_0_I_65 (.A(\DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] ), 
        .B(\DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] ), .C(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] ), .Y(\DWACT_COMP0_E[0] ));
    NOR2A \off_reg_RNIKPQG[0]  (.A(\off_reg[0]_net_1 ), .B(act_ctl_5_8)
        , .Y(\off_time[0] ));
    AND2 un1_counter_0_I_84 (.A(\DWACT_BL_EQUAL_0_E_1[3] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[1] ));
    DFN1C0 cur_pwm (.D(cur_pwm_RNO_2), .CLK(clk_c), .CLR(n_rst_c), .Q(
        primary_5_c));
    XA1B \counter_RNO[12]  (.A(\counter[12]_net_1 ), .B(counter_c11), 
        .C(N_400_0), .Y(counter_n12));
    NOR3C \counter_RNIOLV81[8]  (.A(\counter[7]_net_1 ), .B(counter_c6)
        , .C(\counter[8]_net_1 ), .Y(counter_c8));
    AOI1A un1_counter_0_I_95 (.A(\ACT_LT4_E[3] ), .B(\ACT_LT4_E[6] ), 
        .C(\ACT_LT4_E[10] ), .Y(\DWACT_CMPLE_PO0_DWACT_COMP0_E[0] ));
    OA1A un1_counter_0_I_40 (.A(N_46), .B(N_48), .C(N_47), .Y(N_51));
    XA1B \counter_RNO[1]  (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(N_400_0), .Y(counter_n1));
    DFN1C0 \counter[17]  (.D(counter_n17), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[17]_net_1 ));
    NOR2 un1_counter_2_0_I_129 (.A(\counter[0]_net_1 ), .B(act_ctl_5_4)
        , .Y(N_4));
    DFN1C0 \counter[4]  (.D(counter_n4), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[4]_net_1 ));
    AO1B un1_counter_2_0_I_131 (.A(act_ctl_5_0), .B(\counter[1]_net_1 )
        , .C(N_4), .Y(N_6));
    AND2 un1_counter_0_I_30 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] ));
    OR2A un1_counter_0_I_60 (.A(\counter[23]_net_1 ), .B(
        \off_time[23] ), .Y(N_39));
    DFN1E1C0 \off_reg[11]  (.D(off_div[11]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[11]_net_1 ));
    AND2 un1_counter_0_I_29 (.A(\DWACT_BL_EQUAL_0_E_1[4] ), .B(
        \DWACT_BL_EQUAL_0_E_3[3] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] ));
    NOR2A \off_reg_RNIPUQG[5]  (.A(\off_reg[5]_net_1 ), .B(act_ctl_5_8)
        , .Y(\off_time[5] ));
    DFN1E1C0 \off_reg[22]  (.D(off_div[22]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[22]_net_1 ));
    DFN1C0 \counter[10]  (.D(counter_n10), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[10]_net_1 ));
    NOR2A un1_counter_2_0_I_19 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] ), .B(\counter[31]_net_1 )
        , .Y(\DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] ));
    NOR2A un1_counter_0_I_46 (.A(\off_time[24] ), .B(
        \counter[24]_net_1 ), .Y(\ACT_LT3_E[0] ));
    GND GND_i (.Y(GND));
    DFN1C0 \counter[13]  (.D(counter_n13), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[13]_net_1 ));
    XNOR2 un1_counter_0_I_81 (.A(\counter[16]_net_1 ), .B(
        \off_time[16] ), .Y(\DWACT_BL_EQUAL_0_E_0[1] ));
    NOR2A un1_counter_0_I_90 (.A(\off_time[18] ), .B(
        \counter[18]_net_1 ), .Y(\ACT_LT4_E[5] ));
    XNOR2 un1_counter_0_I_74 (.A(\counter[11]_net_1 ), .B(
        \off_time[11] ), .Y(\DWACT_BL_EQUAL_0_E_1[1] ));
    NOR2B un1_counter_2_0_I_140 (.A(\DWACT_COMP0_E[2] ), .B(
        \DWACT_COMP0_E[1] ), .Y(I_140_5));
    OA1A un1_counter_0_I_36 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .C(N_43), .Y(N_47));
    XNOR2 un1_counter_0_I_66 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\DWACT_BL_EQUAL_0_E[8] ));
    AND3 un1_counter_0_I_17 (.A(\DWACT_BL_EQUAL_0_E_5[0] ), .B(
        \DWACT_BL_EQUAL_0_E_4[1] ), .C(\DWACT_BL_EQUAL_0_E_5[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] ));
    DFN1E1C0 \off_reg[17]  (.D(off_div[17]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[17]_net_1 ));
    AX1C \counter_RNO_0[10]  (.A(\counter[9]_net_1 ), .B(counter_c8), 
        .C(\counter[10]_net_1 ), .Y(counter_n10_tz));
    DFN1C0 \counter[12]  (.D(counter_n12), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[12]_net_1 ));
    OR2A un1_counter_0_I_130 (.A(\off_time[4] ), .B(\counter[4]_net_1 )
        , .Y(N_5));
    NOR2B un1_counter_2_0_I_139 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E[2] )
        , .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ), .Y(
        \DWACT_COMP0_E[2] ));
    NOR2A \off_reg_RNIC21E[27]  (.A(\off_reg[27]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[27] ));
    DFN1C0 \counter[27]  (.D(counter_n27), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[27]_net_1 ));
    OR2A un1_counter_0_I_96 (.A(\off_time[11] ), .B(
        \counter[11]_net_1 ), .Y(N_22));
    NOR2A \off_reg_RNI3MSC[10]  (.A(\off_reg[10]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[10] ));
    NOR2A \off_reg_RNIBUSC[18]  (.A(\off_reg[18]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[18] ));
    AOI1A un1_counter_0_I_49 (.A(\ACT_LT3_E[0] ), .B(\ACT_LT3_E[1] ), 
        .C(\ACT_LT3_E[2] ), .Y(\ACT_LT3_E[3] ));
    NOR2B \counter_RNIOJAC2[14]  (.A(counter_c13), .B(
        \counter[14]_net_1 ), .Y(counter_c14));
    AX1C \counter_RNO_0[20]  (.A(\counter[19]_net_1 ), .B(counter_c18), 
        .C(\counter[20]_net_1 ), .Y(counter_n20_tz));
    DFN1C0 \counter[20]  (.D(counter_n20), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[20]_net_1 ));
    OA1A un1_counter_0_I_101 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .C(N_23), .Y(N_27));
    DFN1E1C0 \off_reg[19]  (.D(off_div[19]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[19]_net_1 ));
    XNOR2 un1_counter_0_I_71 (.A(\counter[10]_net_1 ), .B(
        \off_time[10] ), .Y(\DWACT_BL_EQUAL_0_E_2[0] ));
    OR2A un1_counter_0_I_116 (.A(\off_time[6] ), .B(\counter[6]_net_1 )
        , .Y(N_12));
    AO1C un1_counter_0_I_39 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .C(N_45), .Y(N_50));
    XA1B \counter_RNO[17]  (.A(\counter[17]_net_1 ), .B(counter_c16), 
        .C(N_400_0), .Y(counter_n17));
    XNOR2 un1_counter_0_I_69 (.A(\counter[16]_net_1 ), .B(
        \off_time[16] ), .Y(\DWACT_BL_EQUAL_0_E[6] ));
    XNOR2 un1_counter_0_I_112 (.A(\counter[9]_net_1 ), .B(
        \off_time[9] ), .Y(\DWACT_BL_EQUAL_0_E[4] ));
    OA1A un1_counter_0_I_105 (.A(N_26), .B(N_28), .C(N_27), .Y(N_31));
    DFN1C0 \counter[23]  (.D(counter_n23), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[23]_net_1 ));
    NOR2A \off_reg_RNI6PSC[13]  (.A(\off_reg[13]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[13] ));
    NOR2A \off_reg_RNIATSC[17]  (.A(\off_reg[17]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[17] ));
    NOR2A \off_reg_RNI6QTC[22]  (.A(\off_reg[22]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[22] ));
    XA1B \counter_RNO[29]  (.A(\counter[29]_net_1 ), .B(counter_c28), 
        .C(cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n29));
    DFN1E1C0 \off_reg[25]  (.D(off_div[25]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[25]_net_1 ));
    NOR2B \counter_RNO_0[18]  (.A(counter_c16), .B(\counter[17]_net_1 )
        , .Y(counter_c17));
    DFN1C0 \counter[22]  (.D(counter_n22), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[22]_net_1 ));
    DFN1C0 \counter[15]  (.D(counter_n15), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[15]_net_1 ));
    AO1 un1_counter_0_I_107 (.A(\DWACT_CMPLE_PO0_DWACT_COMP0_E[1] ), 
        .B(\DWACT_CMPLE_PO0_DWACT_COMP0_E[2] ), .C(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] ));
    OR2A un1_counter_0_I_99 (.A(\off_time[14] ), .B(
        \counter[14]_net_1 ), .Y(N_25));
    NOR3C \counter_RNIQGMJ1[10]  (.A(\counter[9]_net_1 ), .B(
        counter_c8), .C(\counter[10]_net_1 ), .Y(counter_c10));
    NOR2A un1_counter_2_0_I_122 (.A(I_20_6), .B(\counter[7]_net_1 ), 
        .Y(N_18));
    AND2 un1_counter_2_0_I_115 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] ));
    XNOR2 un1_counter_0_I_108 (.A(\counter[5]_net_1 ), .B(
        \off_time[5] ), .Y(\DWACT_BL_EQUAL_0_E_0[0] ));
    NOR2B \counter_RNITU195[29]  (.A(counter_c28), .B(
        \counter[29]_net_1 ), .Y(counter_c29));
    AX1C \counter_RNO_0[8]  (.A(\counter[7]_net_1 ), .B(counter_c6), 
        .C(\counter[8]_net_1 ), .Y(counter_n8_tz));
    AX1C \counter_RNO_0[28]  (.A(\counter[27]_net_1 ), .B(counter_c26), 
        .C(\counter[28]_net_1 ), .Y(counter_n28_tz));
    VCC VCC_i (.Y(VCC));
    AO1C un1_counter_0_I_120 (.A(\off_time[6] ), .B(\counter[6]_net_1 )
        , .C(N_14_0), .Y(N_16_0));
    DFN1E1C0 \off_reg[31]  (.D(off_div[31]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[31]_net_1 ));
    XA1B \counter_RNO[14]  (.A(\counter[14]_net_1 ), .B(counter_c13), 
        .C(N_400_0), .Y(counter_n14));
    XNOR2 un1_counter_2_0_I_111 (.A(\counter[7]_net_1 ), .B(I_20_6), 
        .Y(\DWACT_BL_EQUAL_0_E[2] ));
    DFN1E1C0 \off_reg[7]  (.D(off_div[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[7]_net_1 ));
    DFN1C0 \counter[1]  (.D(counter_n1), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[1]_net_1 ));
    XNOR2 un1_counter_0_I_2 (.A(\counter[19]_net_1 ), .B(
        \off_time[19] ), .Y(\DWACT_BL_EQUAL_0_E_5[0] ));
    NOR2A \counter_RNO[26]  (.A(counter_n26_tz), .B(
        cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n26));
    NOR2A un1_counter_0_I_55 (.A(\off_time[19] ), .B(
        \counter[19]_net_1 ), .Y(N_34));
    AO1 un1_counter_0_I_139 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] ), .Y(\DWACT_COMP0_E_0[2] )
        );
    XA1B \counter_RNO[5]  (.A(\counter[5]_net_1 ), .B(counter_c4), .C(
        N_400_0), .Y(counter_n5));
    AO1C un1_counter_0_I_133 (.A(\counter[2]_net_1 ), .B(\off_time[2] )
        , .C(N_2_0), .Y(N_8_0));
    NOR2A \off_reg_RNI7QSC[14]  (.A(\off_reg[14]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[14] ));
    DFN1C0 \counter[25]  (.D(counter_n25), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[25]_net_1 ));
    AND2A un1_counter_0_I_87 (.A(\off_time[16] ), .B(
        \counter[16]_net_1 ), .Y(\ACT_LT4_E[2] ));
    XA1B \counter_RNO[3]  (.A(\counter[3]_net_1 ), .B(counter_c2), .C(
        N_400_0), .Y(counter_n3));
    DFN1E1C0 \off_reg[6]  (.D(off_div[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[6]_net_1 ));
    AND3 un1_counter_0_I_28 (.A(\DWACT_BL_EQUAL_0_E_4[0] ), .B(
        \DWACT_BL_EQUAL_0_E_3[1] ), .C(\DWACT_BL_EQUAL_0_E_4[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] ));
    NOR2A \off_reg_RNI4OTC[20]  (.A(\off_reg[20]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[20] ));
    OR2A un1_counter_0_I_50 (.A(\off_time[26] ), .B(
        \counter[26]_net_1 ), .Y(\ACT_LT3_E[4] ));
    DFN1C0 \counter[5]  (.D(counter_n5), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[5]_net_1 ));
    NOR2A \off_reg_RNIS1RG[8]  (.A(\off_reg[8]_net_1 ), .B(act_ctl_5_8)
        , .Y(\off_time[8] ));
    NOR2A \off_reg_RNIA01E[25]  (.A(\off_reg[25]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[25] ));
    MX2A cur_pwm_RNO (.A(I_140_6), .B(I_140_5), .S(primary_5_c), .Y(
        cur_pwm_RNO_2));
    XNOR2 un1_counter_0_I_4 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(\DWACT_BL_EQUAL_0_E[10] ));
    XNOR2 un1_counter_0_I_23 (.A(\counter[27]_net_1 ), .B(
        \off_time[27] ), .Y(\DWACT_BL_EQUAL_0_E_4[0] ));
    NOR2A \counter_RNO[10]  (.A(counter_n10_tz), .B(
        cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n10));
    AND3 un1_counter_0_I_77 (.A(\DWACT_BL_EQUAL_0_E_2[0] ), .B(
        \DWACT_BL_EQUAL_0_E_1[1] ), .C(\DWACT_BL_EQUAL_0_E_2[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] ));
    XNOR2 un1_counter_0_I_3 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .Y(\DWACT_BL_EQUAL_0_E[11] ));
    XA1B \counter_RNO[21]  (.A(\counter[21]_net_1 ), .B(counter_c20), 
        .C(N_400_0), .Y(counter_n21));
    XNOR2 un1_counter_0_I_6 (.A(\counter[20]_net_1 ), .B(
        \off_time[20] ), .Y(\DWACT_BL_EQUAL_0_E_4[1] ));
    OR2A un1_counter_0_I_56 (.A(\off_time[23] ), .B(
        \counter[23]_net_1 ), .Y(N_35));
    OR2 \off_reg_RNINSQG[3]  (.A(\off_reg[3]_net_1 ), .B(act_ctl_5_8), 
        .Y(\off_time[3] ));
    AX1C \counter_RNO_0[24]  (.A(\counter[23]_net_1 ), .B(counter_c22), 
        .C(\counter[24]_net_1 ), .Y(counter_n24_tz));
    AND3 un1_counter_0_I_15 (.A(\DWACT_BL_EQUAL_0_E_0[6] ), .B(
        \DWACT_BL_EQUAL_0_E_0[7] ), .C(\DWACT_BL_EQUAL_0_E_0[8] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] ));
    NOR2B \counter_RNI0GRP1[11]  (.A(counter_c10), .B(
        \counter[11]_net_1 ), .Y(counter_c11));
    AND2A un1_counter_0_I_48 (.A(\off_time[25] ), .B(
        \counter[25]_net_1 ), .Y(\ACT_LT3_E[2] ));
    NOR2A un1_counter_0_I_129 (.A(\off_time[0] ), .B(
        \counter[0]_net_1 ), .Y(N_4_0));
    XNOR2 un1_counter_0_I_9 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(\DWACT_BL_EQUAL_0_E[12] ));
    AO1 un1_counter_0_I_140 (.A(\DWACT_COMP0_E_0[1] ), .B(
        \DWACT_COMP0_E_0[2] ), .C(\DWACT_COMP0_E[0] ), .Y(I_140_6));
    OR2A un1_counter_0_I_123 (.A(\counter[9]_net_1 ), .B(\off_time[9] )
        , .Y(N_19));
    DFN1C0 \counter[16]  (.D(counter_n16), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[16]_net_1 ));
    OR2A un1_counter_0_I_38 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(N_49));
    XA1B \counter_RNO[25]  (.A(\counter[25]_net_1 ), .B(counter_c24), 
        .C(cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n25));
    XNOR2 un1_counter_0_I_68 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\DWACT_BL_EQUAL_0_E[7] ));
    NOR2A \off_reg_RNI8RSC[15]  (.A(\off_reg[15]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[15] ));
    MX2C cur_pwm_RNIQQ9OA2 (.A(I_140_6), .B(I_140_5), .S(primary_5_c), 
        .Y(N_400_0));
    XNOR2 un1_act_ctl_I_14 (.A(N_5_0), .B(act_ctl_5_4), .Y(I_14_6));
    NOR2B \counter_RNO_0[31]  (.A(\counter[30]_net_1 ), .B(counter_c29)
        , .Y(counter_63_0));
    NOR2B \counter_RNIH3AC[13]  (.A(\counter[13]_net_1 ), .B(
        \counter[14]_net_1 ), .Y(counter_m6_0_a2_2));
    NOR2A \off_reg_RNI5PTC[21]  (.A(\off_reg[21]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[21] ));
    XNOR2 un1_counter_0_I_43 (.A(\counter[25]_net_1 ), .B(
        \off_time[25] ), .Y(\DWACT_BL_EQUAL_0_E_2[1] ));
    XOR2 un1_act_ctl_I_20 (.A(act_ctl_5_4), .B(N_3), .Y(I_20_6));
    AO1C un1_counter_0_I_59 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .C(N_32), .Y(N_38));
    DFN1E1C0 \off_reg[21]  (.D(off_div[21]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[21]_net_1 ));
    AO1C un1_counter_0_I_104 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .C(N_25), .Y(N_30));
    OR2 un1_counter_2_0_I_127 (.A(\counter[1]_net_1 ), .B(act_ctl_5_4), 
        .Y(N_2));
    XNOR2 un1_counter_0_I_10 (.A(\counter[24]_net_1 ), .B(
        \off_time[24] ), .Y(\DWACT_BL_EQUAL_0_E_0[5] ));
    NOR2A un1_counter_0_I_98 (.A(\off_time[10] ), .B(
        \counter[10]_net_1 ), .Y(N_24));
    NOR2A un1_counter_0_I_33 (.A(\off_time[27] ), .B(
        \counter[27]_net_1 ), .Y(N_44));
    OA1 un1_counter_0_I_63 (.A(N_41), .B(N_40), .C(N_39), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] ));
    NOR2A \off_reg_RNI7RTC[23]  (.A(\off_reg[23]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[23] ));
    NOR2A \counter_RNO[6]  (.A(counter_n6_tz), .B(
        cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n6));
    XA1B \counter_RNO[30]  (.A(\counter[30]_net_1 ), .B(counter_c29), 
        .C(cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n30));
    NOR2A \off_reg_RNI6T1E[30]  (.A(\off_reg[30]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[30] ));
    XNOR2 un1_counter_0_I_110 (.A(\counter[8]_net_1 ), .B(
        \off_time[8] ), .Y(\DWACT_BL_EQUAL_0_E_0[3] ));
    DFN1E1C0 \off_reg[27]  (.D(off_div[27]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[27]_net_1 ));
    AND3 un1_counter_0_I_16 (.A(\DWACT_BL_EQUAL_0_E_4[3] ), .B(
        \DWACT_BL_EQUAL_0_E_2[4] ), .C(\DWACT_BL_EQUAL_0_E_0[5] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] ));
    OR2A un1_counter_0_I_93 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\ACT_LT4_E[8] ));
    DFN1E1C0 \off_reg[8]  (.D(off_div[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[8]_net_1 ));
    DFN1C0 \counter[26]  (.D(counter_n26), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[26]_net_1 ));
    XA1B \counter_RNO[23]  (.A(\counter[23]_net_1 ), .B(counter_c22), 
        .C(N_400_0), .Y(counter_n23));
    OA1C un1_counter_2_0_I_137 (.A(\counter[3]_net_1 ), .B(N_11), .C(
        \counter[4]_net_1 ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] ));
    OR2B un1_counter_2_0_I_133 (.A(N_2), .B(\counter[2]_net_1 ), .Y(
        N_8));
    OR2 un1_act_ctl_I_19 (.A(\DWACT_FDEC_E[2] ), .B(\DWACT_FDEC_E[0] ), 
        .Y(N_3));
    DFN1C0 \counter[14]  (.D(counter_n14), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[14]_net_1 ));
    DFN1E1C0 \off_reg[29]  (.D(off_div[29]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[29]_net_1 ));
    AND3 un1_counter_2_0_I_18 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] ));
    DFN1E1C0 \off_reg[1]  (.D(off_div[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[1]_net_1 ));
    NOR2A \counter_RNO[22]  (.A(counter_n22_tz), .B(
        cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n22));
    AO1C un1_counter_0_I_131 (.A(\off_time[1] ), .B(\counter[1]_net_1 )
        , .C(N_4_0), .Y(N_6_0));
    AND2 un1_counter_0_I_19 (.A(\DWACT_BL_EQUAL_0_E[12] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] ));
    XNOR2 un1_counter_0_I_42 (.A(\counter[26]_net_1 ), .B(
        \off_time[26] ), .Y(\DWACT_BL_EQUAL_0_E_3[2] ));
    AO1C un1_counter_0_I_135 (.A(\counter[3]_net_1 ), .B(\off_time[3] )
        , .C(N_5), .Y(N_10));
    NOR2A \off_reg_RNI5OSC[12]  (.A(\off_reg[12]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[12] ));
    DFN1E1C0 \off_reg[10]  (.D(off_div[10]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[10]_net_1 ));
    NOR2A un1_counter_0_I_85 (.A(\off_time[15] ), .B(
        \counter[15]_net_1 ), .Y(\ACT_LT4_E[0] ));
    DFN1C0 \counter[31]  (.D(counter_n31), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[31]_net_1 ));
    OR2A un1_counter_0_I_32 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(N_43));
    OA1A un1_counter_0_I_62 (.A(N_36), .B(N_38), .C(N_37), .Y(N_41));
    OR3A un1_act_ctl_I_13 (.A(act_ctl_5_0), .B(act_ctl_5_0), .C(
        \DWACT_FDEC_E[0] ), .Y(N_5_0));
    OA1 un1_counter_0_I_137 (.A(N_11_0), .B(N_10), .C(N_9), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] ));
    NOR3C \counter_RNIECOM[4]  (.A(\counter[3]_net_1 ), .B(counter_c2), 
        .C(\counter[4]_net_1 ), .Y(counter_c4));
    AO1 un1_counter_0_I_138 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] ));
    NOR2A \off_reg_RNIB11E[26]  (.A(\off_reg[26]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[26] ));
    NOR2A un1_counter_0_I_92 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\ACT_LT4_E[7] ));
    DFN1C0 \counter[24]  (.D(counter_n24), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[24]_net_1 ));
    OR2A un1_counter_0_I_119 (.A(\off_time[9] ), .B(\counter[9]_net_1 )
        , .Y(N_15));
    NOR3 un1_counter_2_0_I_14 (.A(\counter[29]_net_1 ), .B(
        \counter[30]_net_1 ), .C(\counter[28]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] ));
    AND3 un1_counter_2_0_I_78 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ));
    XNOR2 un1_counter_0_I_80 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\DWACT_BL_EQUAL_0_E_1[2] ));
    XNOR2 un1_counter_0_I_5 (.A(\counter[27]_net_1 ), .B(
        \off_time[27] ), .Y(\DWACT_BL_EQUAL_0_E_0[8] ));
    AND3 un1_counter_0_I_113 (.A(\DWACT_BL_EQUAL_0_E_0[0] ), .B(
        \DWACT_BL_EQUAL_0_E[1] ), .C(\DWACT_BL_EQUAL_0_E_0[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] ));
    XNOR2 un1_counter_0_I_24 (.A(\counter[28]_net_1 ), .B(
        \off_time[28] ), .Y(\DWACT_BL_EQUAL_0_E_3[1] ));
    NOR2A \off_reg_RNID31E[28]  (.A(\off_reg[28]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[28] ));
    NOR3C \counter_RNIJHPU[18]  (.A(\counter[16]_net_1 ), .B(
        \counter[18]_net_1 ), .C(counter_m6_0_a2_4), .Y(
        counter_m6_0_a2_6));
    NOR2A \counter_RNO[4]  (.A(counter_n4_tz), .B(
        cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n4));
    AND3 un1_counter_0_I_75 (.A(\DWACT_BL_EQUAL_0_E[6] ), .B(
        \DWACT_BL_EQUAL_0_E[7] ), .C(\DWACT_BL_EQUAL_0_E[8] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] ));
    DFN1E1C0 \off_reg[14]  (.D(off_div[14]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[14]_net_1 ));
    OR2A un1_counter_2_0_I_120 (.A(N_14), .B(\counter[6]_net_1 ), .Y(
        N_16));
    XA1B \counter_RNO[18]  (.A(\counter[18]_net_1 ), .B(counter_c17), 
        .C(N_400_0), .Y(counter_n18));
    NOR3 un1_counter_2_0_I_15 (.A(\counter[26]_net_1 ), .B(
        \counter[27]_net_1 ), .C(\counter[25]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] ));
    OR2A un1_counter_0_I_86 (.A(\off_time[16] ), .B(
        \counter[16]_net_1 ), .Y(\ACT_LT4_E[1] ));
    NOR2A un1_counter_2_0_I_124 (.A(I_23_9), .B(\counter[8]_net_1 ), 
        .Y(N_20));
    OA1A un1_counter_0_I_58 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .C(N_33), .Y(N_37));
    OA1A un1_counter_0_I_121 (.A(\counter[8]_net_1 ), .B(\off_time[8] )
        , .C(N_13_0), .Y(N_17_0));
    AND2 un1_counter_2_0_I_20 (.A(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] ), .B(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] ), .Y(
        \DWACT_COMP0_E[1] ));
    AX1C \counter_RNO_0[26]  (.A(\counter[25]_net_1 ), .B(counter_c24), 
        .C(\counter[26]_net_1 ), .Y(counter_n26_tz));
    XA1B \counter_RNO[27]  (.A(\counter[27]_net_1 ), .B(counter_c26), 
        .C(cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n27));
    OA1A un1_counter_0_I_125 (.A(N_16_0), .B(N_18_0), .C(N_17_0), .Y(
        N_21_0));
    NOR3C \counter_RNIHKDN1[11]  (.A(counter_m6_0_a2_2), .B(
        counter_m6_0_a2_1), .C(counter_m6_0_a2_6), .Y(
        counter_m6_0_a2_7));
    AX1C \counter_RNO_0[6]  (.A(\counter[5]_net_1 ), .B(counter_c4), 
        .C(\counter[6]_net_1 ), .Y(counter_n6_tz));
    NOR2B \counter_RNIDRKO2[16]  (.A(counter_c15), .B(
        \counter[16]_net_1 ), .Y(counter_c16));
    XNOR2 un1_counter_0_I_70 (.A(\counter[15]_net_1 ), .B(
        \off_time[15] ), .Y(\DWACT_BL_EQUAL_0_E[5] ));
    OA1 un1_counter_0_I_106 (.A(N_31), .B(N_30), .C(N_29), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] ));
    DFN1E1C0 \off_reg[18]  (.D(off_div[18]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[18]_net_1 ));
    AO1C un1_counter_0_I_102 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .C(N_22), .Y(N_28));
    OR2A un1_counter_2_0_I_117 (.A(\counter[7]_net_1 ), .B(I_20_6), .Y(
        N_13));
    NOR3B un1_counter_2_0_I_113 (.A(\DWACT_BL_EQUAL_0_E[2] ), .B(
        \DWACT_BL_EQUAL_0_E[0] ), .C(\counter[6]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ));
    XNOR2 un1_counter_0_I_44 (.A(\counter[24]_net_1 ), .B(
        \off_time[24] ), .Y(\DWACT_BL_EQUAL_0_E_3[0] ));
    OR2A un1_counter_0_I_53 (.A(\off_time[20] ), .B(
        \counter[20]_net_1 ), .Y(N_32));
    OR2A un1_counter_0_I_127 (.A(\off_time[1] ), .B(\counter[1]_net_1 )
        , .Y(N_2_0));
    OR2A un1_counter_0_I_34 (.A(\off_time[31] ), .B(
        \counter[31]_net_1 ), .Y(N_45));
    OR2A un1_counter_0_I_128 (.A(\counter[2]_net_1 ), .B(\off_time[2] )
        , .Y(N_3_0));
    NOR3C \counter_RNIVTKD[2]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .C(\counter[2]_net_1 ), .Y(counter_c2));
    OR2A un1_counter_0_I_89 (.A(\off_time[17] ), .B(
        \counter[17]_net_1 ), .Y(\ACT_LT4_E[4] ));
    AO1 un1_counter_0_I_64 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] ));
    DFN1E1C0 \off_reg[16]  (.D(off_div[16]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[16]_net_1 ));
    AND3 un1_counter_0_I_76 (.A(\DWACT_BL_EQUAL_0_E_2[3] ), .B(
        \DWACT_BL_EQUAL_0_E_0[4] ), .C(\DWACT_BL_EQUAL_0_E[5] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] ));
    NOR2A \off_reg_RNIE41E[29]  (.A(\off_reg[29]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[29] ));
    XNOR2 un1_counter_0_I_1 (.A(\counter[23]_net_1 ), .B(
        \off_time[23] ), .Y(\DWACT_BL_EQUAL_0_E_2[4] ));
    DFN1E1C0 \off_reg[30]  (.D(off_div[30]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[30]_net_1 ));
    NOR3 un1_counter_2_0_I_75 (.A(\counter[17]_net_1 ), .B(
        \counter[18]_net_1 ), .C(\counter[16]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] ));
    NOR2A \counter_RNO[24]  (.A(counter_n24_tz), .B(
        cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n24));
    DFN1C0 \counter[7]  (.D(counter_n7), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[7]_net_1 ));
    AOI1A un1_counter_0_I_94 (.A(\ACT_LT4_E[7] ), .B(\ACT_LT4_E[8] ), 
        .C(\ACT_LT4_E[5] ), .Y(\ACT_LT4_E[10] ));
    DFN1C0 \counter[30]  (.D(counter_n30), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[30]_net_1 ));
    OA1 un1_counter_0_I_41 (.A(N_51), .B(N_50), .C(N_49), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] ));
    NOR2A \off_reg_RNI8STC[24]  (.A(\off_reg[24]_net_1 ), .B(
        act_ctl_5_6), .Y(\off_time[24] ));
    AND3 un1_counter_0_I_18 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] ));
    NOR3C \counter_RNIQEAH3[19]  (.A(\counter[19]_net_1 ), .B(
        counter_c18), .C(\counter[20]_net_1 ), .Y(counter_c20));
    OR2A un1_counter_0_I_31 (.A(\off_time[28] ), .B(
        \counter[28]_net_1 ), .Y(N_42));
    XNOR2 un1_counter_2_0_I_108 (.A(\counter[5]_net_1 ), .B(I_14_6), 
        .Y(\DWACT_BL_EQUAL_0_E[0] ));
    AO1C un1_counter_0_I_61 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .C(N_35), .Y(N_40));
    NOR2 \counter_RNO[0]  (.A(\counter[0]_net_1 ), .B(
        cur_pwm_RNIQQ9OA2_0_net_1), .Y(\counter_RNO_2[0] ));
    XNOR2 un1_counter_0_I_79 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\DWACT_BL_EQUAL_0_E_1[3] ));
    NOR2B \counter_RNIFH562[13]  (.A(counter_c12), .B(
        \counter[13]_net_1 ), .Y(counter_c13));
    DFN1E1C0 \off_reg[3]  (.D(off_div[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[3]_net_1 ));
    NOR2A \off_reg_RNIT2RG[9]  (.A(\off_reg[9]_net_1 ), .B(act_ctl_5_8)
        , .Y(\off_time[9] ));
    DFN1E1C0 \off_reg[0]  (.D(off_div[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[0]_net_1 ));
    OR3 un1_act_ctl_I_18 (.A(act_ctl_5_0), .B(act_ctl_5_i), .C(
        act_ctl_5_1), .Y(\DWACT_FDEC_E[2] ));
    OA1B un1_counter_2_0_I_126 (.A(N_20), .B(N_21), .C(
        \counter[9]_net_1 ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ));
    OR2A un1_counter_0_I_134 (.A(\counter[4]_net_1 ), .B(\off_time[4] )
        , .Y(N_9));
    XNOR2 un1_counter_0_I_13 (.A(\counter[28]_net_1 ), .B(
        \off_time[28] ), .Y(\DWACT_BL_EQUAL_0_E[9] ));
    NOR2A un1_counter_0_I_91 (.A(\ACT_LT4_E[4] ), .B(\ACT_LT4_E[5] ), 
        .Y(\ACT_LT4_E[6] ));
    AOI1A un1_counter_0_I_52 (.A(\ACT_LT3_E[3] ), .B(\ACT_LT3_E[4] ), 
        .C(\ACT_LT3_E[5] ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] ));
    NOR3C \counter_RNIR6FI[10]  (.A(\counter[15]_net_1 ), .B(
        \counter[10]_net_1 ), .C(\counter[17]_net_1 ), .Y(
        counter_m6_0_a2_4));
    NOR3C \counter_RNI9IMT3[22]  (.A(\counter[21]_net_1 ), .B(
        counter_c20), .C(\counter[22]_net_1 ), .Y(counter_c22));
    NOR2A \counter_RNO[20]  (.A(counter_n20_tz), .B(
        cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n20));
    DFN1E1C0 \off_reg[13]  (.D(off_div[13]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[13]_net_1 ));
    XNOR2 un1_counter_0_I_27 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(\DWACT_BL_EQUAL_0_E_1[4] ));
    XNOR2 un1_counter_0_I_111 (.A(\counter[7]_net_1 ), .B(
        \off_time[7] ), .Y(\DWACT_BL_EQUAL_0_E_0[2] ));
    OR2A un1_counter_2_0_I_136 (.A(N_6), .B(N_8), .Y(N_11));
    OR2 \off_reg_RNIMRQG[2]  (.A(\off_reg[2]_net_1 ), .B(act_ctl_5_8), 
        .Y(\off_time[2] ));
    AND2 un1_counter_0_I_115 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] ));
    DFN1E1C0 \off_reg[4]  (.D(off_div[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg), .Q(\off_reg[4]_net_1 ));
    XNOR2 un1_counter_2_0_I_110 (.A(\counter[8]_net_1 ), .B(I_23_9), 
        .Y(\DWACT_BL_EQUAL_0_E[3] ));
    XNOR2 un1_counter_0_I_8 (.A(\counter[25]_net_1 ), .B(
        \off_time[25] ), .Y(\DWACT_BL_EQUAL_0_E_0[6] ));
    DFN1E1C0 \off_reg[20]  (.D(off_div[20]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[20]_net_1 ));
    NOR2A \counter_RNO[2]  (.A(counter_n2_tz), .B(
        cur_pwm_RNIQQ9OA2_0_net_1), .Y(counter_n2));
    DFN1C0 \counter[9]  (.D(counter_n9), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[9]_net_1 ));
    NOR3 un1_counter_2_0_I_16 (.A(\counter[24]_net_1 ), .B(
        \counter[23]_net_1 ), .C(\counter[22]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] ));
    NOR2A un1_counter_2_0_I_114 (.A(\DWACT_BL_EQUAL_0_E[3] ), .B(
        \counter[9]_net_1 ), .Y(\DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ));
    OR2A un1_counter_0_I_117 (.A(\counter[7]_net_1 ), .B(\off_time[7] )
        , .Y(N_13_0));
    XA1B \counter_RNO[19]  (.A(\counter[19]_net_1 ), .B(counter_c18), 
        .C(N_400_0), .Y(counter_n19));
    AO1C un1_counter_0_I_124 (.A(\counter[8]_net_1 ), .B(\off_time[8] )
        , .C(N_15), .Y(N_20_0));
    NOR2A un1_counter_0_I_118 (.A(\off_time[5] ), .B(
        \counter[5]_net_1 ), .Y(N_14_0));
    XNOR2 un1_counter_0_I_12 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .Y(\DWACT_BL_EQUAL_0_E_5[2] ));
    AO1 un1_counter_2_0_I_138 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] )
        , .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] ));
    XA1B \counter_RNO[9]  (.A(\counter[9]_net_1 ), .B(counter_c8), .C(
        N_400_0), .Y(counter_n9));
    DFN1E1C0 \off_reg[12]  (.D(off_div[12]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[12]_net_1 ));
    AOI1A un1_counter_0_I_88 (.A(\ACT_LT4_E[0] ), .B(\ACT_LT4_E[1] ), 
        .C(\ACT_LT4_E[2] ), .Y(\ACT_LT4_E[3] ));
    OR2A un1_counter_0_I_47 (.A(\off_time[25] ), .B(
        \counter[25]_net_1 ), .Y(\ACT_LT3_E[1] ));
    NOR3C \counter_RNI1VRV[5]  (.A(\counter[5]_net_1 ), .B(counter_c4), 
        .C(\counter[6]_net_1 ), .Y(counter_c6));
    DFN1C0 \counter[8]  (.D(counter_n8), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[8]_net_1 ));
    OR2A un1_counter_0_I_54 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .Y(N_33));
    AO1C un1_counter_0_I_37 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .C(N_42), .Y(N_48));
    NOR3C \counter_RNIELR25[27]  (.A(\counter[27]_net_1 ), .B(
        counter_c26), .C(\counter[28]_net_1 ), .Y(counter_c28));
    XNOR2 un1_counter_0_I_7 (.A(\counter[26]_net_1 ), .B(
        \off_time[26] ), .Y(\DWACT_BL_EQUAL_0_E_0[7] ));
    XNOR2 un1_counter_0_I_67 (.A(\counter[14]_net_1 ), .B(
        \off_time[14] ), .Y(\DWACT_BL_EQUAL_0_E_0[4] ));
    DFN1C0 \counter[18]  (.D(counter_n18), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[18]_net_1 ));
    AO1C un1_counter_0_I_100 (.A(\off_time[11] ), .B(
        \counter[11]_net_1 ), .C(N_24), .Y(N_26));
    OR2 \off_reg_RNILQQG[1]  (.A(\off_reg[1]_net_1 ), .B(act_ctl_5_8), 
        .Y(\off_time[1] ));
    DFN1E1C0 \off_reg[24]  (.D(off_div[24]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[24]_net_1 ));
    AND3 un1_counter_0_I_83 (.A(\DWACT_BL_EQUAL_0_E_1[0] ), .B(
        \DWACT_BL_EQUAL_0_E_0[1] ), .C(\DWACT_BL_EQUAL_0_E_1[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] ));
    XA1B \counter_RNO[16]  (.A(\counter[16]_net_1 ), .B(counter_c15), 
        .C(N_400_0), .Y(counter_n16));
    DFN1C0 \counter[0]  (.D(\counter_RNO_2[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\counter[0]_net_1 ));
    NOR3 un1_counter_2_0_I_76 (.A(\counter[15]_net_1 ), .B(
        \counter[14]_net_1 ), .C(\counter[13]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] ));
    OR2A un1_counter_0_I_97 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .Y(N_23));
    
endmodule


module spi_clk_11s_2(
       sck_fb_c,
       n_rst_c,
       clk_c
    );
output sck_fb_c;
input  n_rst_c;
input  clk_c;

    wire N_8, \counter[1]_net_1 , \counter[0]_net_1 , N_6, 
        \counter[3]_net_1 , \DWACT_FINC_E[0] , cur_clk5_5, cur_clk5_3, 
        \counter[6]_net_1 , cur_clk5_4, cur_clk5_1, \counter[7]_net_1 , 
        \counter[8]_net_1 , \counter[4]_net_1 , \counter[5]_net_1 , 
        \counter[2]_net_1 , cur_clk_RNO_2, \counter_3[1] , I_5_2, 
        \counter_3[0] , \counter_3[3] , I_9_2, I_7_2, I_12_3, I_14_5, 
        I_17_3, I_20_5, I_23_7, N_2, \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[3] , N_3, N_4, \DWACT_FINC_E[1] , N_5, N_7, GND, 
        VCC;
    
    NOR2B un3_counter_I_6 (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(N_8));
    AND3 un3_counter_I_19 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\counter[6]_net_1 ), .Y(N_3));
    XOR2 un3_counter_I_20 (.A(N_3), .B(\counter[7]_net_1 ), .Y(I_20_5));
    DFN1C0 \counter[2]  (.D(I_7_2), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[2]_net_1 ));
    DFN1C0 \counter[7]  (.D(I_20_5), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[7]_net_1 ));
    AND3 un3_counter_I_13 (.A(\DWACT_FINC_E[0] ), .B(
        \counter[3]_net_1 ), .C(\counter[4]_net_1 ), .Y(N_5));
    AOI1 \counter_RNO[0]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(
        \counter[0]_net_1 ), .Y(\counter_3[0] ));
    DFN1C0 \counter[6]  (.D(I_17_3), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[6]_net_1 ));
    NOR3A \counter_RNI2ELU[8]  (.A(cur_clk5_1), .B(\counter[7]_net_1 ), 
        .C(\counter[8]_net_1 ), .Y(cur_clk5_4));
    VCC VCC_i (.Y(VCC));
    XOR2 un3_counter_I_12 (.A(N_6), .B(\counter[4]_net_1 ), .Y(I_12_3));
    DFN1C0 \counter[8]  (.D(I_23_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[8]_net_1 ));
    XOR2 un3_counter_I_23 (.A(N_2), .B(\counter[8]_net_1 ), .Y(I_23_7));
    AOI1B \counter_RNO[1]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(I_5_2), 
        .Y(\counter_3[1] ));
    AND3 un3_counter_I_22 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\DWACT_FINC_E[3] ), .Y(N_2));
    XOR2 un3_counter_I_7 (.A(N_8), .B(\counter[2]_net_1 ), .Y(I_7_2));
    NOR2B un3_counter_I_11 (.A(\counter[3]_net_1 ), .B(
        \DWACT_FINC_E[0] ), .Y(N_6));
    AND3 un3_counter_I_16 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[1] )
        , .C(\counter[5]_net_1 ), .Y(N_4));
    DFN1C0 \counter[4]  (.D(I_12_3), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[4]_net_1 ));
    XOR2 un3_counter_I_17 (.A(N_4), .B(\counter[6]_net_1 ), .Y(I_17_3));
    DFN1C0 \counter[5]  (.D(I_14_5), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[5]_net_1 ));
    AND3 un3_counter_I_8 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(N_7));
    GND GND_i (.Y(GND));
    AX1C cur_clk_RNO (.A(cur_clk5_4), .B(cur_clk5_5), .C(sck_fb_c), .Y(
        cur_clk_RNO_2));
    AOI1B \counter_RNO[3]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(I_9_2), 
        .Y(\counter_3[3] ));
    AND2 un3_counter_I_21 (.A(\counter[6]_net_1 ), .B(
        \counter[7]_net_1 ), .Y(\DWACT_FINC_E[3] ));
    DFN1C0 \counter[1]  (.D(\counter_3[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[1]_net_1 ));
    DFN1C0 \counter[3]  (.D(\counter_3[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[3]_net_1 ));
    NOR3B \counter_RNIQ5LU[6]  (.A(\counter[1]_net_1 ), .B(cur_clk5_3), 
        .C(\counter[6]_net_1 ), .Y(cur_clk5_5));
    AND2 un3_counter_I_15 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(\DWACT_FINC_E[1] ));
    XOR2 un3_counter_I_9 (.A(N_7), .B(\counter[3]_net_1 ), .Y(I_9_2));
    DFN1C0 cur_clk (.D(cur_clk_RNO_2), .CLK(clk_c), .CLR(n_rst_c), .Q(
        sck_fb_c));
    NOR2A \counter_RNITIAF[4]  (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(cur_clk5_3));
    XOR2 un3_counter_I_14 (.A(N_5), .B(\counter[5]_net_1 ), .Y(I_14_5));
    NOR2 \counter_RNITIAF[2]  (.A(\counter[5]_net_1 ), .B(
        \counter[2]_net_1 ), .Y(cur_clk5_1));
    XOR2 un3_counter_I_5 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .Y(I_5_2));
    AND3 un3_counter_I_10 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(
        \DWACT_FINC_E[0] ));
    DFN1C0 \counter[0]  (.D(\counter_3[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[0]_net_1 ));
    AND3 un3_counter_I_18 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .C(\counter[5]_net_1 ), .Y(
        \DWACT_FINC_E[2] ));
    
endmodule


module PID_controller_Z4(
       choose_0_0,
       LED_12_0,
       LED_12_2,
       LED_12_3,
       LED_12_5,
       LED_15_0,
       LED_15_2,
       LED_15_3,
       LED_15_5,
       LED_c_0,
       LED_c_2,
       LED_c_5,
       choose,
       LED_FB_0,
       LED_FB_2,
       LED_FB_5,
       LED_33_0,
       LED_33_2,
       LED_33_5,
       LED_5_0,
       LED_5_3,
       LED_5_5,
       LED_5_6,
       primary_5_c,
       act_ctl_5_4,
       act_ctl_5_8,
       act_ctl_5_6,
       act_ctl_5_7,
       act_ctl_5_0,
       act_ctl_5_1,
       act_ctl_5_i,
       N_45,
       din_5_c,
       cs_i_1_i,
       sck_fb_c,
       clk_c,
       n_rst_c
    );
input  choose_0_0;
input  LED_12_0;
input  LED_12_2;
input  LED_12_3;
input  LED_12_5;
input  LED_15_0;
input  LED_15_2;
input  LED_15_3;
input  LED_15_5;
output LED_c_0;
output LED_c_2;
output LED_c_5;
input  [2:0] choose;
input  LED_FB_0;
input  LED_FB_2;
input  LED_FB_5;
input  LED_33_0;
input  LED_33_2;
input  LED_33_5;
output LED_5_0;
output LED_5_3;
output LED_5_5;
output LED_5_6;
output primary_5_c;
input  act_ctl_5_4;
input  act_ctl_5_8;
input  act_ctl_5_6;
input  act_ctl_5_7;
input  act_ctl_5_0;
input  act_ctl_5_1;
input  act_ctl_5_i;
output N_45;
input  din_5_c;
output cs_i_1_i;
output sck_fb_c;
input  clk_c;
input  n_rst_c;

    wire \state[0] , \state[1] , pwm_chg, sig_prev, sig_old_i_0, 
        avg_done, N_46_1, vd_rdy, sum_rdy, deriv_enable, calc_avg, 
        calc_int, pwm_enable, sum_enable, calc_error, avg_enable, 
        int_enable, pwm_chg_0, avg_enable_0, avg_enable_1, \cur_vd[0] , 
        \cur_vd[1] , \cur_vd[2] , \cur_vd[3] , \cur_vd[4] , 
        \cur_vd[5] , \cur_vd[6] , \cur_vd[7] , \cur_vd[8] , 
        \cur_vd[9] , \cur_vd[10] , \cur_vd[11] , \avg_new[0] , 
        \avg_new[1] , \avg_new[2] , \avg_new[3] , \avg_new[4] , 
        \avg_new[5] , \avg_new[6] , \avg_new[7] , \avg_new[8] , 
        \avg_new[9] , \avg_new[10] , \avg_new[11] , \avg_old[0] , 
        \avg_old[1] , \avg_old[2] , \avg_old[3] , \avg_old[4] , 
        \avg_old[5] , \avg_old[6] , \avg_old[7] , \avg_old[8] , 
        \avg_old[9] , \avg_old[10] , \avg_old[11] , \cur_error[0] , 
        \cur_error[1] , \cur_error[2] , \cur_error[3] , \cur_error[4] , 
        \cur_error[5] , \cur_error[6] , \cur_error[7] , \cur_error[8] , 
        \cur_error[9] , \cur_error[10] , \cur_error[11] , 
        \cur_error[12] , \LED_5_i[5] , \LED_5[0] , \LED_5[2] , 
        \LED_5[3] , \LED_5[5] , \average[2] , \average[3] , 
        \average[4] , \average[5] , \average[6] , \sr_old[0] , 
        \sr_old[1] , \sr_old[2] , \sr_old[3] , \sr_old[4] , 
        \sr_old[5] , \sr_old[6] , \sr_old[7] , \sr_old[8] , 
        \sr_old[9] , \sr_old[10] , \sr_old[11] , \sr_old[12] , 
        \sr_new[0] , \sr_new[1] , \sr_new[2] , \sr_new[3] , 
        \sr_new[4] , \sr_new[5] , \sr_new[6] , \sr_new[7] , 
        \sr_new[8] , \sr_new[9] , \sr_new[10] , \sr_new[11] , 
        \sr_new[12] , \sr_prev[0] , \sr_prev[1] , \sr_prev[2] , 
        \sr_prev[3] , \sr_prev[4] , \sr_prev[5] , \sr_prev[6] , 
        \sr_prev[7] , \sr_prev[8] , \sr_prev[9] , \sr_prev[10] , 
        \sr_prev[11] , \sr_prev[12] , \sr_new_0[12] , \sr_new_1[12] , 
        \integral[6] , \integral[7] , \integral[8] , \integral[9] , 
        \integral[10] , \integral[11] , \integral[12] , \integral[13] , 
        \integral[14] , \integral[15] , \integral[16] , \integral[17] , 
        \integral[18] , \integral[19] , \integral[20] , \integral[21] , 
        \integral[22] , \integral[23] , \integral[24] , \integral[25] , 
        \integral_i[24] , \integral_i[25] , \integral_0[25] , 
        \integral_1[25] , \derivative[12] , \sum[39] , \sum[14] , 
        \sum[19] , \sum[20] , \sum[22] , \sum[13] , \sum[17] , 
        \sum[18] , \sum[23] , \sum[21] , \sum[16] , \sum[15] , 
        \sum[12] , \sum[11] , \sum[6] , \sum[10] , \sum[9] , \sum[5] , 
        \sum[8] , \sum[7] , \sum[4] , \sum[2] , \sum[1] , \sum[0] , 
        \sum[3] , \sum_0[39] , \sum_1[39] , \sum_2[39] , vd_done, 
        \off_div[0] , \off_div[1] , \off_div[2] , \off_div[3] , 
        \off_div[4] , \off_div[5] , \off_div[6] , \off_div[7] , 
        \off_div[8] , \off_div[9] , \off_div[10] , \off_div[11] , 
        \off_div[12] , \off_div[13] , \off_div[14] , \off_div[15] , 
        \off_div[16] , \off_div[17] , \off_div[18] , \off_div[19] , 
        \off_div[20] , \off_div[21] , \off_div[22] , \off_div[23] , 
        \off_div[24] , \off_div[25] , \off_div[26] , \off_div[27] , 
        \off_div[28] , \off_div[29] , \off_div[30] , \off_div[31] , 
        GND, VCC;
    
    pwm_ctl_400s_32s_13s_0_1_2_4 PWM_CTL (.sum_8(\sum[8] ), .sum_39(
        \sum[39] ), .sum_10(\sum[10] ), .sum_11(\sum[11] ), .sum_12(
        \sum[12] ), .sum_13(\sum[13] ), .sum_14(\sum[14] ), .sum_16(
        \sum[16] ), .sum_17(\sum[17] ), .sum_18(\sum[18] ), .sum_19(
        \sum[19] ), .sum_20(\sum[20] ), .sum_21(\sum[21] ), .sum_22(
        \sum[22] ), .sum_23(\sum[23] ), .sum_15(\sum[15] ), .sum_9(
        \sum[9] ), .sum_0_d0(\sum[0] ), .sum_2_d0(\sum[2] ), .sum_1_d0(
        \sum[1] ), .sum_7(\sum[7] ), .sum_6(\sum[6] ), .sum_4(\sum[4] )
        , .sum_3(\sum[3] ), .sum_5(\sum[5] ), .LED_33_0(LED_33_0), 
        .LED_33_2(LED_33_2), .LED_33_5(LED_33_5), .LED_FB_0(LED_FB_0), 
        .LED_FB_2(LED_FB_2), .LED_FB_5(LED_FB_5), .LED_5_0(\LED_5[0] ), 
        .LED_5_2(\LED_5[2] ), .LED_5_3(\LED_5[3] ), .LED_5_5(
        \LED_5[5] ), .choose({choose[2], choose[1], choose[0]}), 
        .LED_c_0(LED_c_0), .LED_c_2(LED_c_2), .LED_c_5(LED_c_5), 
        .LED_15_0(LED_15_0), .LED_15_2(LED_15_2), .LED_15_3(LED_15_3), 
        .LED_15_5(LED_15_5), .LED_12_0(LED_12_0), .LED_12_2(LED_12_2), 
        .LED_12_3(LED_12_3), .LED_12_5(LED_12_5), .choose_0_0(
        choose_0_0), .off_div({\off_div[31] , \off_div[30] , 
        \off_div[29] , \off_div[28] , \off_div[27] , \off_div[26] , 
        \off_div[25] , \off_div[24] , \off_div[23] , \off_div[22] , 
        \off_div[21] , \off_div[20] , \off_div[19] , \off_div[18] , 
        \off_div[17] , \off_div[16] , \off_div[15] , \off_div[14] , 
        \off_div[13] , \off_div[12] , \off_div[11] , \off_div[10] , 
        \off_div[9] , \off_div[8] , \off_div[7] , \off_div[6] , 
        \off_div[5] , \off_div[4] , \off_div[3] , \off_div[2] , 
        \off_div[1] , \off_div[0] }), .sum_1_0(\sum_1[39] ), .sum_0_0(
        \sum_0[39] ), .sum_2_0(\sum_2[39] ), .state({\state[1] , 
        \state[0] }), .n_rst_c(n_rst_c), .clk_c(clk_c), .N_45(N_45), 
        .pwm_enable(pwm_enable));
    integral_calc_13s_4_2 AVG_CALC (.avg_old({\avg_old[11] , 
        \avg_old[10] , \avg_old[9] , \avg_old[8] , \avg_old[7] , 
        \avg_old[6] , \avg_old[5] , \avg_old[4] , \avg_old[3] , 
        \avg_old[2] , \avg_old[1] , \avg_old[0] }), .avg_new({
        \avg_new[11] , \avg_new[10] , \avg_new[9] , \avg_new[8] , 
        \avg_new[7] , \avg_new[6] , \avg_new[5] , \avg_new[4] , 
        \avg_new[3] , \avg_new[2] , \avg_new[1] , \avg_new[0] }), 
        .LED_5({LED_5_6, LED_5_5, \LED_5[5] , LED_5_3, \LED_5[3] , 
        \LED_5[2] , LED_5_0, \LED_5[0] }), .average({\average[6] , 
        \average[5] , \average[4] , \average[3] , \average[2] }), 
        .LED_5_i_0(\LED_5_i[5] ), .calc_avg(calc_avg), .avg_done(
        avg_done), .n_rst_c(n_rst_c), .clk_c(clk_c));
    error_sr_13s_5s_2 AVGSR (.cur_vd({\cur_vd[11] , \cur_vd[10] , 
        \cur_vd[9] , \cur_vd[8] , \cur_vd[7] , \cur_vd[6] , 
        \cur_vd[5] , \cur_vd[4] , \cur_vd[3] , \cur_vd[2] , 
        \cur_vd[1] , \cur_vd[0] }), .avg_new({\avg_new[11] , 
        \avg_new[10] , \avg_new[9] , \avg_new[8] , \avg_new[7] , 
        \avg_new[6] , \avg_new[5] , \avg_new[4] , \avg_new[3] , 
        \avg_new[2] , \avg_new[1] , \avg_new[0] }), .avg_old({
        \avg_old[11] , \avg_old[10] , \avg_old[9] , \avg_old[8] , 
        \avg_old[7] , \avg_old[6] , \avg_old[5] , \avg_old[4] , 
        \avg_old[3] , \avg_old[2] , \avg_old[1] , \avg_old[0] }), 
        .avg_enable_1(avg_enable_1), .avg_enable_0(avg_enable_0), 
        .avg_enable(avg_enable), .n_rst_c(n_rst_c), .clk_c(clk_c));
    error_sr_13s_64s_2 INTSR (.sr_old({\sr_old[12] , \sr_old[11] , 
        \sr_old[10] , \sr_old[9] , \sr_old[8] , \sr_old[7] , 
        \sr_old[6] , \sr_old[5] , \sr_old[4] , \sr_old[3] , 
        \sr_old[2] , \sr_old[1] , \sr_old[0] }), .sr_new({\sr_new[12] , 
        \sr_new[11] , \sr_new[10] , \sr_new[9] , \sr_new[8] , 
        \sr_new[7] , \sr_new[6] , \sr_new[5] , \sr_new[4] , 
        \sr_new[3] , \sr_new[2] , \sr_new[1] , \sr_new[0] }), 
        .cur_error({\cur_error[12] , \cur_error[11] , \cur_error[10] , 
        \cur_error[9] , \cur_error[8] , \cur_error[7] , \cur_error[6] , 
        \cur_error[5] , \cur_error[4] , \cur_error[3] , \cur_error[2] , 
        \cur_error[1] , \cur_error[0] }), .sr_prev({\sr_prev[12] , 
        \sr_prev[11] , \sr_prev[10] , \sr_prev[9] , \sr_prev[8] , 
        \sr_prev[7] , \sr_prev[6] , \sr_prev[5] , \sr_prev[4] , 
        \sr_prev[3] , \sr_prev[2] , \sr_prev[1] , \sr_prev[0] }), 
        .sr_new_0_0(\sr_new_0[12] ), .sr_new_1_0(\sr_new_1[12] ), 
        .int_enable(int_enable), .n_rst_c(n_rst_c), .clk_c(clk_c));
    controller_Z1_4_2 CONTROLLER (.state_0_0(\state[0] ), .state_0_d0(
        \state[1] ), .pwm_chg(pwm_chg), .sig_prev(sig_prev), 
        .sig_old_i_0(sig_old_i_0), .avg_done(avg_done), .N_46_1(N_46_1)
        , .vd_rdy(vd_rdy), .sum_rdy(sum_rdy), .deriv_enable(
        deriv_enable), .calc_avg(calc_avg), .calc_int(calc_int), 
        .pwm_enable(pwm_enable), .sum_enable(sum_enable), .calc_error(
        calc_error), .avg_enable(avg_enable), .int_enable(int_enable), 
        .pwm_chg_0(pwm_chg_0), .avg_enable_0(avg_enable_0), .n_rst_c(
        n_rst_c), .clk_c(clk_c), .avg_enable_1(avg_enable_1));
    sig_gen_6 FM_CYCLE (.primary_5_c(primary_5_c), .n_rst_c(n_rst_c), 
        .clk_c(clk_c), .sig_old_i_0(sig_old_i_0), .sig_prev(sig_prev));
    pid_sum_13s_4_2 SUM (.integral_i({\integral_i[25] , 
        \integral_i[24] }), .integral({\integral[25] , \integral[24] , 
        \integral[23] , \integral[22] , \integral[21] , \integral[20] , 
        \integral[19] , \integral[18] , \integral[17] , \integral[16] , 
        \integral[15] , \integral[14] , \integral[13] , \integral[12] , 
        \integral[11] , \integral[10] , \integral[9] , \integral[8] , 
        \integral[7] , \integral[6] }), .sr_new({\sr_new[12] , 
        \sr_new[11] , \sr_new[10] , \sr_new[9] , \sr_new[8] , 
        \sr_new[7] , \sr_new[6] , \sr_new[5] , \sr_new[4] , 
        \sr_new[3] , \sr_new[2] , \sr_new[1] , \sr_new[0] }), 
        .integral_1_0(\integral_1[25] ), .sr_new_1_0(\sr_new_1[12] ), 
        .sr_new_0_0(\sr_new_0[12] ), .derivative_0(\derivative[12] ), 
        .integral_0_0(\integral_0[25] ), .sum_39(\sum[39] ), .sum_14(
        \sum[14] ), .sum_19(\sum[19] ), .sum_20(\sum[20] ), .sum_22(
        \sum[22] ), .sum_13(\sum[13] ), .sum_17(\sum[17] ), .sum_18(
        \sum[18] ), .sum_23(\sum[23] ), .sum_21(\sum[21] ), .sum_16(
        \sum[16] ), .sum_15(\sum[15] ), .sum_12(\sum[12] ), .sum_11(
        \sum[11] ), .sum_6(\sum[6] ), .sum_10(\sum[10] ), .sum_9(
        \sum[9] ), .sum_5(\sum[5] ), .sum_8(\sum[8] ), .sum_7(\sum[7] )
        , .sum_4(\sum[4] ), .sum_2_d0(\sum[2] ), .sum_1_d0(\sum[1] ), 
        .sum_0_d0(\sum[0] ), .sum_3(\sum[3] ), .sum_0_0(\sum_0[39] ), 
        .sum_1_0(\sum_1[39] ), .sum_2_0(\sum_2[39] ), .sum_enable(
        sum_enable), .sum_rdy(sum_rdy), .n_rst_c(n_rst_c), .clk_c(
        clk_c));
    sig_gen_5 VD_SIG (.vd_done(vd_done), .n_rst_c(n_rst_c), .clk_c(
        clk_c), .vd_rdy(vd_rdy));
    spi_rx_12s_2 SPI (.cur_vd({\cur_vd[11] , \cur_vd[10] , \cur_vd[9] , 
        \cur_vd[8] , \cur_vd[7] , \cur_vd[6] , \cur_vd[5] , 
        \cur_vd[4] , \cur_vd[3] , \cur_vd[2] , \cur_vd[1] , 
        \cur_vd[0] }), .vd_done(vd_done), .cs_i_1_i(cs_i_1_i), 
        .sck_fb_c(sck_fb_c), .n_rst_c(n_rst_c), .din_5_c(din_5_c));
    integral_calc_13s_0_4_2 INTCALC (.sr_new({\sr_new[12] , 
        \sr_new[11] , \sr_new[10] , \sr_new[9] , \sr_new[8] , 
        \sr_new[7] , \sr_new[6] , \sr_new[5] , \sr_new[4] , 
        \sr_new[3] , \sr_new[2] , \sr_new[1] , \sr_new[0] }), .sr_old({
        \sr_old[12] , \sr_old[11] , \sr_old[10] , \sr_old[9] , 
        \sr_old[8] , \sr_old[7] , \sr_old[6] , \sr_old[5] , 
        \sr_old[4] , \sr_old[3] , \sr_old[2] , \sr_old[1] , 
        \sr_old[0] }), .sr_new_0_0(\sr_new_0[12] ), .sr_new_1_0(
        \sr_new_1[12] ), .integral({\integral[25] , \integral[24] , 
        \integral[23] , \integral[22] , \integral[21] , \integral[20] , 
        \integral[19] , \integral[18] , \integral[17] , \integral[16] , 
        \integral[15] , \integral[14] , \integral[13] , \integral[12] , 
        \integral[11] , \integral[10] , \integral[9] , \integral[8] , 
        \integral[7] , \integral[6] }), .integral_i({\integral_i[25] , 
        \integral_i[24] }), .integral_0_0(\integral_0[25] ), 
        .integral_1_0(\integral_1[25] ), .calc_int(calc_int), .N_46_1(
        N_46_1), .n_rst_c(n_rst_c), .clk_c(clk_c));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    error_calc_13s_12s_4_2 EC (.cur_error({\cur_error[12] , 
        \cur_error[11] , \cur_error[10] , \cur_error[9] , 
        \cur_error[8] , \cur_error[7] , \cur_error[6] , \cur_error[5] , 
        \cur_error[4] , \cur_error[3] , \cur_error[2] , \cur_error[1] , 
        \cur_error[0] }), .LED_5_i_0(\LED_5_i[5] ), .LED_5({LED_5_6, 
        LED_5_5, \LED_5[5] , LED_5_3, \LED_5[3] , \LED_5[2] , LED_5_0, 
        \LED_5[0] }), .average({\average[6] , \average[5] , 
        \average[4] , \average[3] , \average[2] }), .calc_error(
        calc_error), .n_rst_c(n_rst_c), .clk_c(clk_c));
    derivative_calc_13s_4_2 DCALC (.derivative_0(\derivative[12] ), 
        .sr_prev({\sr_prev[12] , \sr_prev[11] , \sr_prev[10] , 
        \sr_prev[9] , \sr_prev[8] , \sr_prev[7] , \sr_prev[6] , 
        \sr_prev[5] , \sr_prev[4] , \sr_prev[3] , \sr_prev[2] , 
        \sr_prev[1] , \sr_prev[0] }), .sr_new({\sr_new[11] , 
        \sr_new[10] , \sr_new[9] , \sr_new[8] , \sr_new[7] , 
        \sr_new[6] , \sr_new[5] , \sr_new[4] , \sr_new[3] , 
        \sr_new[2] , \sr_new[1] , \sr_new[0] }), .sr_new_0_0(
        \sr_new_0[12] ), .deriv_enable(deriv_enable), .n_rst_c(n_rst_c)
        , .clk_c(clk_c));
    pwm_tx_400s_32s_13s_10_222s_45s PWM_TX (.off_div({\off_div[31] , 
        \off_div[30] , \off_div[29] , \off_div[28] , \off_div[27] , 
        \off_div[26] , \off_div[25] , \off_div[24] , \off_div[23] , 
        \off_div[22] , \off_div[21] , \off_div[20] , \off_div[19] , 
        \off_div[18] , \off_div[17] , \off_div[16] , \off_div[15] , 
        \off_div[14] , \off_div[13] , \off_div[12] , \off_div[11] , 
        \off_div[10] , \off_div[9] , \off_div[8] , \off_div[7] , 
        \off_div[6] , \off_div[5] , \off_div[4] , \off_div[3] , 
        \off_div[2] , \off_div[1] , \off_div[0] }), .act_ctl_5_i(
        act_ctl_5_i), .act_ctl_5_1(act_ctl_5_1), .act_ctl_5_0(
        act_ctl_5_0), .pwm_chg_0(pwm_chg_0), .pwm_chg(pwm_chg), 
        .n_rst_c(n_rst_c), .clk_c(clk_c), .act_ctl_5_7(act_ctl_5_7), 
        .act_ctl_5_6(act_ctl_5_6), .act_ctl_5_8(act_ctl_5_8), 
        .act_ctl_5_4(act_ctl_5_4), .primary_5_c(primary_5_c));
    spi_clk_11s_2 SPICLK (.sck_fb_c(sck_fb_c), .n_rst_c(n_rst_c), 
        .clk_c(clk_c));
    
endmodule


module pwm_ctl_200s_32s_13s_0_1_2_1(
       sum_8,
       sum_39,
       sum_12,
       sum_14,
       sum_15,
       sum_16,
       sum_17,
       sum_18,
       sum_21,
       sum_22,
       sum_23,
       sum_9,
       sum_10,
       sum_19,
       sum_11,
       sum_20,
       sum_13,
       sum_1_d0,
       sum_0_d0,
       sum_2_d0,
       sum_7,
       sum_6,
       sum_3,
       sum_5,
       sum_4,
       sum_0_0,
       off_div,
       sum_1_0,
       sum_2_0,
       state,
       n_rst_c,
       clk_c,
       pwm_enable
    );
input  sum_8;
input  sum_39;
input  sum_12;
input  sum_14;
input  sum_15;
input  sum_16;
input  sum_17;
input  sum_18;
input  sum_21;
input  sum_22;
input  sum_23;
input  sum_9;
input  sum_10;
input  sum_19;
input  sum_11;
input  sum_20;
input  sum_13;
input  sum_1_d0;
input  sum_0_d0;
input  sum_2_d0;
input  sum_7;
input  sum_6;
input  sum_3;
input  sum_5;
input  sum_4;
input  sum_0_0;
output [31:0] off_div;
input  sum_1_0;
input  sum_2_0;
output [1:0] state;
input  n_rst_c;
input  clk_c;
input  pwm_enable;

    wire un1_state_2_0, un5lt31, next_off_div_2_sqmuxa_10, 
        \state_d_0[2] , N_16, \DWACT_FINC_E[4] , N_13, 
        \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , ADD_32x32_fast_I321_Y_0, 
        ADD_32x32_fast_I258_Y_3, N610, N625, ADD_32x32_fast_I258_Y_2, 
        N482, ADD_32x32_fast_I258_Y_0, N551, ADD_32x32_fast_I320_Y_0, 
        ADD_32x32_fast_I313_Y_0, ADD_32x32_fast_I259_Y_3, N627, N612, 
        ADD_32x32_fast_I259_Y_2, N553, N546, ADD_32x32_fast_I259_Y_1, 
        N484, N481, ADD_32x32_fast_I259_Y_0, 
        ADD_32x32_fast_I258_un1_Y_0, N626, ADD_32x32_fast_I319_Y_0, 
        ADD_32x32_fast_I318_Y_0, ADD_32x32_fast_I317_Y_0, 
        ADD_32x32_fast_I316_Y_0, ADD_32x32_fast_I315_Y_0, 
        ADD_32x32_fast_I314_Y_0, ADD_32x32_fast_I266_Y_0, N641, 
        ADD_32x32_fast_I261_Y_2, N616, N631, ADD_32x32_fast_I261_Y_1, 
        N488, N557, ADD_32x32_fast_I260_Y_2, N629, N614, 
        ADD_32x32_fast_I260_Y_1, N555, N548, ADD_32x32_fast_I260_Y_0, 
        N486, ADD_32x32_fast_I312_Y_0, ADD_32x32_fast_I304_Y_0, 
        \sum_adj[22]_net_1 , ADD_32x32_fast_I259_un1_Y_0, N628, 
        ADD_32x32_fast_I262_Y_1, N618, N633, ADD_32x32_fast_I262_Y_0, 
        N559, ADD_32x32_fast_I311_Y_0, ADD_32x32_fast_I310_Y_0, 
        ADD_32x32_fast_I309_Y_0, ADD_32x32_fast_I266_un1_Y_0, N642, 
        ADD_32x32_fast_I264_Y_1, N622, N637, ADD_32x32_fast_I264_Y_0, 
        N563, ADD_32x32_fast_I265_Y_0, N558, N565, 
        ADD_32x32_fast_I263_Y_1, N620, N635, ADD_32x32_fast_I263_Y_0, 
        N561, ADD_32x32_fast_I306_Y_0, ADD_32x32_fast_I307_Y_0, 
        ADD_32x32_fast_I308_Y_0, ADD_32x32_fast_I302_Y_0, 
        \un1_sum_adj[12] , ADD_32x32_fast_I303_Y_0, \un1_sum_adj[13] , 
        ADD_32x32_fast_I260_un1_Y_0, N630, ADD_32x32_fast_I261_un1_Y_0, 
        N632, ADD_32x32_fast_I301_Y_0, \sum_adj[19]_net_1 , 
        ADD_32x32_fast_I262_un1_Y_0, N634, ADD_32x32_fast_I269_Y_0, 
        N647, ADD_32x32_fast_I270_Y_0, N649, ADD_32x32_fast_I299_Y_0, 
        \un1_sum_adj[9] , ADD_32x32_fast_I300_Y_0, \un1_sum_adj[10] , 
        ADD_32x32_fast_I298_Y_0, \un1_sum_adj[8] , 
        ADD_32x32_fast_I264_un1_Y_0, N638, ADD_32x32_fast_I265_un1_Y_0, 
        N624, N640, ADD_32x32_fast_I263_un1_Y_0, N636, 
        ADD_32x32_fast_I296_Y_0, \un1_sum_adj[6] , 
        ADD_32x32_fast_I271_Y_0, ADD_32x32_fast_I271_un1_Y_0, 
        ADD_32x32_fast_I272_Y_0, ADD_32x32_fast_I272_un1_Y_0, 
        ADD_32x32_fast_I273_Y_0, ADD_32x32_fast_I273_un1_Y_0, N639, 
        ADD_32x32_fast_I295_Y_0, \sum_adj[13]_net_1 , 
        ADD_32x32_fast_I294_Y_0, \un1_sum_adj[4] , 
        ADD_32x32_fast_I293_Y_0, \sum_adj[11]_net_1 , N538, N654, N590, 
        N598, \sum_adj_RNISG3M[8]_net_1 , N586, N594, N601, 
        ADD_32x32_fast_I292_Y_0, \un1_sum_adj[2] , 
        next_off_div_2_sqmuxa_8, next_off_div_2_sqmuxa_7, 
        next_off_div16, next_off_div_2_sqmuxa_2, 
        next_off_div_2_sqmuxa_1, next_off_div_2_sqmuxa_5, 
        next_off_div_2_sqmuxa_4, ADD_32x32_fast_I291_Y_0, 
        \sum_adj[9]_net_1 , un5lto20_2, un5lto20_1, 
        ADD_32x32_fast_I155_Y_0, un5lto14_2, un5lto14_1, 
        un1_off_divlto31_22, un1_off_divlto31_15, un1_off_divlto31_14, 
        un1_off_divlto31_20, un1_off_divlto31_21, un1_off_divlto31_13, 
        un1_off_divlto31_12, un1_off_divlto31_17, un1_off_divlto31_10, 
        un1_off_divlto31_9, un1_off_divlt31, un1_off_divlto31_0, 
        un5lto9, un1_off_divlto31_8, un1_off_divlto31_6, 
        un1_off_divlto31_4, un1_off_divlto31_2, un5lto7_1, N483, N552, 
        \un1_off_div_1[0] , N749, N781, \un1_off_div_1[17] , 
        I238_un1_Y, N757, N793, N769, I230_un1_Y, I268_un1_Y, N646, 
        N661, N761, N799, N765, N657, \un1_off_div_1[18] , I236_un1_Y, 
        \un1_off_div_1[7] , \un1_sum_adj[7] , N759, N796, I270_un1_Y, 
        N650, N599, \un1_off_div_1[3] , \un1_off_div_1[5] , 
        \un1_off_div_1[19] , N755, N790, N485, N489, 
        \un1_off_div_1[10] , I269_un1_Y, N648, N663, 
        \un1_off_div_1[20] , \un1_off_div_1[15] , \un1_sum_adj[15] , 
        N751, N784, N779, N655, un5lt16, N753, N787, I265_un1_Y, N802, 
        N763, I224_un1_Y, I267_un1_Y, N644, N659, N767, I228_un1_Y, 
        un5lt9, un5lto4, un5lt4, \nsum_adj_5[8] , I_23_0, 
        \nsum_adj_5[12] , I_35, \nsum_adj_5[14] , I_40, 
        \nsum_adj_5[15] , I_43, \nsum_adj_5[16] , I_46, 
        \nsum_adj_5[17] , I_49, \nsum_adj_5[18] , I_53, 
        \nsum_adj_5[21] , I_62, \nsum_adj_5[22] , I_65, 
        \nsum_adj_5[23] , I_70, state_176_d, \nsum_adj_5[9] , I_26, 
        N_311_i, \nsum_adj_5[10] , I_28, N643, N556, 
        \next_off_div[29] , \state_d[2] , \next_off_div[24] , 
        \next_off_div[22] , \nsum_adj_5[19] , I_56, \nsum_adj_5[11] , 
        I_32, \state_RNIURLQM_0[1]_net_1 , un5lt14, \nsum_adj_5[20] , 
        I_59, \nsum_adj_5[13] , I_37, N493, \next_off_div[30] , 
        \next_off_div[16] , \state_ns[0] , \next_off_div[6] , 
        \next_off_div[8] , \next_off_div[11] , \next_off_div[13] , 
        \next_off_div[14] , N383, N521, N411, N524, N401, N405, N404, 
        N534, N386, N390, N389, N535, N387, N536, N537, 
        \sum_adj[8]_net_1 , N525, N589, N528, N529, N595, N531, N530, 
        N596, N407, N416, N417, N422, N425, N426, N428, N429, N508, 
        N509, N510, N511, N513, N420, N573, N512, N574, N582, N517, 
        I184_un1_Y, N581, \sum_adj[23]_net_1 , \sum_adj[21]_net_1 , 
        \sum_adj[16]_net_1 , \next_off_div[15] , next_off_div_1_sqmuxa, 
        \sum_adj[10]_net_1 , I150_un1_Y, N645, N432, N506, N507, 
        \next_off_div[20] , \sum_adj[20]_net_1 , N566, N419, N597, 
        N533, N532, \next_off_div[2] , \sum_adj[14]_net_1 , 
        \sum_adj[15]_net_1 , N523, \next_off_div[10] , N526, N398, 
        N527, N399, N584, N519, N587, N522, N588, N591, N514, N502, 
        N498, N572, N571, N564, N503, N499, N494, N495, N496, N497, 
        N560, N567, N568, N491, \next_off_div[12] , \next_off_div[28] , 
        N576, N592, N575, N583, \next_off_div[3] , 
        next_off_div_0_sqmuxa, \next_off_div[5] , \next_off_div[19] , 
        \sum_adj[17]_net_1 , \sum_adj[18]_net_1 , N518, N520, N410, 
        N516, N413, N515, N579, N593, N580, N395, \next_off_div[9] , 
        \next_off_div[1] , \next_off_div[26] , N562, N651, I247_un1_Y, 
        \next_off_div[18] , \next_off_div[7] , \next_off_div[23] , 
        N500, N492, N501, N505, N435, N504, I196_un1_Y, N585, N578, 
        N577, N570, N569, N393, N392, \next_off_div[25] , N487, N490, 
        \next_off_div[21] , \next_off_div[27] , I190_un1_Y, 
        \next_off_div[17] , \sum_adj[12]_net_1 , N653, I204_un1_Y, 
        \next_off_div[4] , \next_off_div[31] , \next_off_div[0] , 
        I249_un1_Y, N_2, \DWACT_FINC_E[29] , \DWACT_FINC_E[13] , 
        \DWACT_FINC_E[33] , \DWACT_FINC_E[34] , \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[5] , \DWACT_FINC_E[15] , N_3, \DWACT_FINC_E[28] , 
        \DWACT_FINC_E[16] , N_4, N_5, \DWACT_FINC_E[14] , N_6, 
        \DWACT_FINC_E[9] , \DWACT_FINC_E[12] , N_7, \DWACT_FINC_E[10] , 
        \DWACT_FINC_E[0] , N_8, \DWACT_FINC_E[11] , N_9, N_10, N_11, 
        \DWACT_FINC_E[8] , N_12, N_14, N_15, \DWACT_FINC_E[3] , N_17, 
        GND, VCC;
    
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I59_Y (.A(N435), .B(N432), 
        .Y(N505));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_2 (.A(N482), .B(
        ADD_32x32_fast_I258_Y_0), .C(N551), .Y(ADD_32x32_fast_I258_Y_2)
        );
    DFN1C0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(state[0]));
    DFN1E0C0 \off_div[29]  (.D(\next_off_div[29] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[29]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y_0 (.A(N555), .B(N563), 
        .Y(ADD_32x32_fast_I264_Y_0));
    DFN1E0C0 \off_div[26]  (.D(\next_off_div[26] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[26]));
    XNOR2 un1_nsum_adj_I_43 (.A(sum_15), .B(N_10), .Y(I_43));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I247_Y (.A(I247_un1_Y), .B(
        N651), .Y(N796));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I108_Y (.A(N496), .B(N492), 
        .Y(N557));
    AND3 un1_nsum_adj_I_48 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[11] ), .Y(N_8));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I47_Y (.A(off_div[23]), .B(
        off_div[22]), .C(sum_0_0), .Y(N493));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I3_P0N (.A(sum_2_0), .B(
        \sum_adj[11]_net_1 ), .C(off_div[3]), .Y(N393));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I165_Y (.A(N489), .B(N493), 
        .C(N562), .Y(N620));
    DFN1E0C0 \off_div[31]  (.D(\next_off_div[31] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[31]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I149_Y (.A(N537), .B(N533), 
        .Y(N598));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I135_Y (.A(N519), .B(N523), 
        .Y(N584));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I147_Y (.A(N535), .B(N531), 
        .Y(N596));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I121_Y (.A(N505), .B(N509), 
        .Y(N570));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I272_Y_0 (.A(
        ADD_32x32_fast_I272_un1_Y_0), .B(N638), .C(N637), .Y(
        ADD_32x32_fast_I272_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I173_Y (.A(N562), .B(N570), 
        .Y(N628));
    MX2 \sum_adj_RNO[9]  (.A(sum_9), .B(I_26), .S(sum_2_0), .Y(
        \nsum_adj_5[9] ));
    XA1 \off_div_RNO[22]  (.A(N767), .B(ADD_32x32_fast_I312_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[22] ));
    DFN1E1C0 \sum_adj[23]  (.D(\nsum_adj_5[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[23]_net_1 ));
    NOR3 un1_nsum_adj_I_41 (.A(sum_13), .B(sum_12), .C(sum_14), .Y(
        \DWACT_FINC_E[9] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I203_Y (.A(N594), .B(N601), 
        .C(N593), .Y(N659));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I155_Y (.A(N483), .B(
        ADD_32x32_fast_I155_Y_0), .C(N552), .Y(N610));
    NOR2B un1_nsum_adj_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_13));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I86_Y (.A(N389), .B(N393), .C(
        N392), .Y(N532));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I200_Y (.A(N597), .B(N590), 
        .C(N589), .Y(N655));
    XNOR2 un1_nsum_adj_I_37 (.A(sum_13), .B(N_12), .Y(I_37));
    MX2 \sum_adj_RNO[15]  (.A(sum_15), .B(I_43), .S(sum_2_0), .Y(
        \nsum_adj_5[15] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I315_Y_0 (.A(off_div[25]), 
        .B(sum_39), .Y(ADD_32x32_fast_I315_Y_0));
    NOR3 un1_nsum_adj_I_10 (.A(sum_1_d0), .B(sum_0_d0), .C(sum_2_d0), 
        .Y(\DWACT_FINC_E[0] ));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I84_Y (.A(N392), .B(
        off_div[4]), .C(\un1_sum_adj[4] ), .Y(N530));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I130_Y (.A(N518), .B(N515), 
        .C(N514), .Y(N579));
    NOR2B \off_div_RNIO1HT[19]  (.A(off_div[20]), .B(off_div[19]), .Y(
        un5lto20_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I266_Y (.A(
        ADD_32x32_fast_I266_un1_Y_0), .B(N657), .C(
        ADD_32x32_fast_I266_Y_0), .Y(N765));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I118_Y (.A(N506), .B(N503), 
        .C(N502), .Y(N567));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I273_un1_Y_0 (.A(N590), .B(
        N598), .C(\sum_adj_RNISG3M[8]_net_1 ), .Y(
        ADD_32x32_fast_I273_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I69_Y (.A(N420), .B(N417), 
        .Y(N515));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I262_Y_0 (.A(N551), .B(N559), 
        .Y(ADD_32x32_fast_I262_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I202_Y (.A(N592), .B(N599), 
        .C(N591), .Y(N657));
    MX2 \sum_adj_RNO[16]  (.A(sum_16), .B(I_46), .S(sum_2_0), .Y(
        \nsum_adj_5[16] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I309_Y_0 (.A(off_div[19]), 
        .B(sum_39), .Y(ADD_32x32_fast_I309_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I184_un1_Y (.A(N581), .B(
        N574), .Y(I184_un1_Y));
    NOR3A \off_div_RNIF44R1[22]  (.A(next_off_div_2_sqmuxa_4), .B(
        off_div[22]), .C(off_div[23]), .Y(next_off_div_2_sqmuxa_7));
    OR2B \off_div_RNIEOSF[5]  (.A(off_div[5]), .B(un5lto4), .Y(
        un1_off_divlt31));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I5_P0N (.A(sum_1_0), .B(
        \sum_adj[13]_net_1 ), .C(off_div[5]), .Y(N399));
    MX2 \off_div_RNO[3]  (.A(next_off_div_0_sqmuxa), .B(
        \un1_off_div_1[3] ), .S(\state_d_0[2] ), .Y(\next_off_div[3] ));
    OA1 \off_div_RNI5FSF[1]  (.A(off_div[1]), .B(off_div[0]), .C(
        off_div[2]), .Y(un5lt4));
    XNOR2 un1_nsum_adj_I_70 (.A(sum_23), .B(N_2), .Y(I_70));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I76_Y (.A(N404), .B(
        off_div[8]), .C(\un1_sum_adj[8] ), .Y(N522));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I4_G0N (.A(\un1_sum_adj[4] )
        , .B(off_div[4]), .Y(N395));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I1_P0N (.A(sum_1_0), .B(
        \sum_adj[9]_net_1 ), .C(off_div[1]), .Y(N387));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I13_G0N (.A(
        \un1_sum_adj[13] ), .B(off_div[13]), .Y(N422));
    DFN1E0C0 \off_div[15]  (.D(\next_off_div[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[15]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I150_Y (.A(I150_un1_Y), .B(
        N534), .Y(N599));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I144_Y (.A(N532), .B(N529), 
        .C(N528), .Y(N593));
    XOR2 \sum_adj_RNISG3M[8]  (.A(\sum_adj[8]_net_1 ), .B(sum_2_0), .Y(
        \sum_adj_RNISG3M[8]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I74_Y (.A(N407), .B(N411), .C(
        N410), .Y(N520));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I50_Y (.A(off_div[21]), .B(
        off_div[20]), .C(sum_0_0), .Y(N496));
    DFN1E0C0 \off_div[13]  (.D(\next_off_div[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[13]));
    XNOR2 un1_nsum_adj_I_62 (.A(sum_21), .B(N_4), .Y(I_62));
    MX2 \sum_adj_RNO[20]  (.A(sum_20), .B(I_59), .S(sum_2_0), .Y(
        \nsum_adj_5[20] ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I293_Y_0 (.A(sum_1_0), .B(
        \sum_adj[11]_net_1 ), .C(off_div[3]), .Y(
        ADD_32x32_fast_I293_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I272_un1_Y_0 (.A(N538), .B(
        N654), .Y(ADD_32x32_fast_I272_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I265_un1_Y (.A(
        ADD_32x32_fast_I265_un1_Y_0), .B(N802), .Y(I265_un1_Y));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I319_Y_0 (.A(off_div[29]), 
        .B(sum_39), .Y(ADD_32x32_fast_I319_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I265_Y_0 (.A(N558), .B(N565), 
        .C(N557), .Y(ADD_32x32_fast_I265_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I179_Y (.A(N576), .B(N568), 
        .Y(N634));
    XA1 \off_div_RNO[24]  (.A(N763), .B(ADD_32x32_fast_I314_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[24] ));
    XNOR2 un1_nsum_adj_I_35 (.A(sum_12), .B(N_13), .Y(I_35));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I309_Y (.A(I270_un1_Y), .B(
        ADD_32x32_fast_I270_Y_0), .C(ADD_32x32_fast_I309_Y_0), .Y(
        \un1_off_div_1[19] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I177_Y (.A(N566), .B(N574), 
        .Y(N632));
    XOR2 \sum_adj_RNI5RNQ[10]  (.A(\sum_adj[10]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[2] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I51_Y (.A(off_div[21]), .B(
        off_div[20]), .C(sum_0_0), .Y(N497));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I308_Y_0 (.A(off_div[18]), 
        .B(sum_39), .Y(ADD_32x32_fast_I308_Y_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I2_P0N (.A(\un1_sum_adj[2] ), 
        .B(off_div[2]), .Y(N390));
    DFN1E0P0 \off_div[7]  (.D(\next_off_div[7] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[7]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I196_Y (.A(I196_un1_Y), .B(
        N585), .Y(N651));
    AND3 un1_nsum_adj_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[6] ));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I268_Y (.A(I230_un1_Y), .B(
        N629), .C(I268_un1_Y), .Y(N769));
    DFN1E0C0 \off_div[9]  (.D(\next_off_div[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[9]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I37_Y (.A(off_div[28]), .B(
        off_div[27]), .C(sum_0_0), .Y(N483));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_1 (.A(N484), .B(N481), 
        .C(ADD_32x32_fast_I259_Y_0), .Y(ADD_32x32_fast_I259_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I186_Y (.A(N583), .B(N576), 
        .C(N575), .Y(N641));
    XOR2 \sum_adj_RNI9VNQ[14]  (.A(\sum_adj[14]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[6] ));
    DFN1E0C0 \off_div[11]  (.D(\next_off_div[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[11]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I145_Y (.A(N533), .B(N529), 
        .Y(N594));
    NOR2A un1_nsum_adj_I_63 (.A(\DWACT_FINC_E[15] ), .B(sum_21), .Y(
        \DWACT_FINC_E[16] ));
    DFN1E1C0 \sum_adj[18]  (.D(\nsum_adj_5[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[18]_net_1 ));
    MX2 un1_off_div_1_0_0_ADD_32x32_fast_I92_Y (.A(sum_1_0), .B(
        off_div[0]), .S(\sum_adj[8]_net_1 ), .Y(N538));
    AND3 un1_nsum_adj_I_68 (.A(\DWACT_FINC_E[34] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[29] ));
    XA1 \off_div_RNO[13]  (.A(N787), .B(ADD_32x32_fast_I303_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[13] ));
    NOR2 \off_div_RNI5I1K[7]  (.A(off_div[11]), .B(off_div[7]), .Y(
        un1_off_divlto31_10));
    OR2 \off_div_RNITEJA[9]  (.A(off_div[9]), .B(off_div[8]), .Y(
        un5lto9));
    MX2 \sum_adj_RNO[21]  (.A(sum_21), .B(I_62), .S(sum_2_0), .Y(
        \nsum_adj_5[21] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I318_Y_0 (.A(off_div[28]), 
        .B(sum_39), .Y(ADD_32x32_fast_I318_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I191_Y (.A(N588), .B(N580), 
        .Y(N646));
    MX2 \sum_adj_RNO[22]  (.A(sum_22), .B(I_65), .S(sum_2_0), .Y(
        \nsum_adj_5[22] ));
    MX2 \off_div_RNO[15]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[15] ), .S(\state_d_0[2] ), .Y(
        \next_off_div[15] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y (.A(
        ADD_32x32_fast_I258_un1_Y_0), .B(N781), .C(
        ADD_32x32_fast_I258_Y_3), .Y(N749));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I14_P0N (.A(sum_0_0), .B(
        \sum_adj[22]_net_1 ), .C(off_div[14]), .Y(N426));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I122_Y (.A(N510), .B(N507), 
        .C(N506), .Y(N571));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I89_Y (.A(N390), .B(N387), 
        .Y(N535));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I262_Y_1 (.A(N618), .B(N633), 
        .C(ADD_32x32_fast_I262_Y_0), .Y(ADD_32x32_fast_I262_Y_1));
    AND2 un1_nsum_adj_I_44 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[9] ), .Y(\DWACT_FINC_E[10] ));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I265_Y (.A(I224_un1_Y), .B(
        ADD_32x32_fast_I265_Y_0), .C(I265_un1_Y), .Y(N763));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I181_Y (.A(N570), .B(N578), 
        .Y(N636));
    AND3 un1_nsum_adj_I_61 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[15] ), .Y(N_4));
    NOR2 un1_nsum_adj_I_47 (.A(sum_15), .B(sum_16), .Y(
        \DWACT_FINC_E[11] ));
    DFN1E1C0 \sum_adj[9]  (.D(\nsum_adj_5[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[9]_net_1 ));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I60_Y (.A(N428), .B(sum_1_0), 
        .C(off_div[16]), .Y(N506));
    NOR3A \off_div_RNIJ51R1[18]  (.A(un1_off_divlto31_6), .B(
        off_div[18]), .C(off_div[20]), .Y(un1_off_divlto31_14));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I307_Y (.A(I238_un1_Y), .B(
        ADD_32x32_fast_I272_Y_0), .C(ADD_32x32_fast_I307_Y_0), .Y(
        \un1_off_div_1[17] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I174_Y (.A(N571), .B(N564), 
        .C(N563), .Y(N629));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I140_Y (.A(N528), .B(N525), 
        .C(N524), .Y(N589));
    DFN1E1C0 \sum_adj[11]  (.D(\nsum_adj_5[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[11]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y_1 (.A(N620), .B(N635), 
        .C(ADD_32x32_fast_I263_Y_0), .Y(ADD_32x32_fast_I263_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I246_Y (.A(N650), .B(N599), 
        .C(N649), .Y(N793));
    XA1 \off_div_RNO[27]  (.A(N757), .B(ADD_32x32_fast_I317_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[27] ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I291_Y_0 (.A(sum_1_0), .B(
        \sum_adj[9]_net_1 ), .C(off_div[1]), .Y(
        ADD_32x32_fast_I291_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I249_un1_Y (.A(N590), .B(
        N598), .C(\sum_adj_RNISG3M[8]_net_1 ), .Y(I249_un1_Y));
    NOR3B un1_nsum_adj_I_36 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .C(sum_12), .Y(N_12));
    DFN1E0C0 \off_div[25]  (.D(\next_off_div[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[25]));
    XA1 \off_div_RNO[1]  (.A(N538), .B(ADD_32x32_fast_I291_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[1] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I61_Y (.A(N432), .B(N429), 
        .Y(N507));
    DFN1E1C0 \sum_adj[22]  (.D(\nsum_adj_5[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[22]_net_1 ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I79_Y (.A(off_div[6]), .B(
        \un1_sum_adj[6] ), .C(N405), .Y(N525));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I150_un1_Y (.A(N535), .B(
        N538), .Y(I150_un1_Y));
    DFN1E0C0 \off_div[23]  (.D(\next_off_div[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[23]));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I304_Y_0 (.A(sum_1_0), .B(
        \sum_adj[22]_net_1 ), .C(off_div[14]), .Y(
        ADD_32x32_fast_I304_Y_0));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I298_Y_0 (.A(off_div[8]), .B(
        \un1_sum_adj[8] ), .Y(ADD_32x32_fast_I298_Y_0));
    XA1 \off_div_RNO[9]  (.A(N799), .B(ADD_32x32_fast_I299_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[9] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y_1 (.A(N622), .B(N637), 
        .C(ADD_32x32_fast_I264_Y_0), .Y(ADD_32x32_fast_I264_Y_1));
    GND GND_i (.Y(GND));
    DFN1E1C0 \sum_adj[14]  (.D(\nsum_adj_5[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[14]_net_1 ));
    NOR3B \off_div_RNIVAL0G[22]  (.A(next_off_div_2_sqmuxa_8), .B(
        next_off_div_2_sqmuxa_7), .C(next_off_div16), .Y(
        next_off_div_2_sqmuxa_10));
    NOR2 \off_div_RNIP3IT[24]  (.A(off_div[25]), .B(off_div[24]), .Y(
        next_off_div_2_sqmuxa_2));
    OA1 \off_div_RNI2KFD4[15]  (.A(un5lt14), .B(un5lto14_2), .C(
        off_div[15]), .Y(un5lt16));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I138_Y (.A(N526), .B(N523), 
        .C(N522), .Y(N587));
    NOR2 \off_div_RNIO2IT[22]  (.A(off_div[26]), .B(off_div[22]), .Y(
        un1_off_divlto31_2));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y (.A(
        ADD_32x32_fast_I259_un1_Y_0), .B(N784), .C(
        ADD_32x32_fast_I259_Y_3), .Y(N751));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I43_Y (.A(off_div[25]), .B(
        off_div[24]), .C(sum_0_0), .Y(N489));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I123_Y (.A(N511), .B(N507), 
        .Y(N572));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I175_Y (.A(N564), .B(N572), 
        .Y(N630));
    NOR3B un1_nsum_adj_I_45 (.A(\DWACT_FINC_E[10] ), .B(
        \DWACT_FINC_E[6] ), .C(sum_15), .Y(N_9));
    OA1 \off_div_RNICICA1[1]  (.A(un5lto4), .B(un5lt4), .C(un5lto7_1), 
        .Y(un5lt9));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I106_Y (.A(N494), .B(N490), 
        .Y(N555));
    MX2 \sum_adj_RNO[10]  (.A(sum_10), .B(I_28), .S(sum_1_0), .Y(
        \nsum_adj_5[10] ));
    NOR3A \off_div_RNIJ9GD1[6]  (.A(un1_off_divlto31_0), .B(off_div[6])
        , .C(un5lto9), .Y(un1_off_divlto31_17));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I11_G0N (.A(sum_1_0), .B(
        \sum_adj[19]_net_1 ), .C(off_div[11]), .Y(N416));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I314_Y_0 (.A(off_div[24]), 
        .B(sum_39), .Y(ADD_32x32_fast_I314_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I271_un1_Y_0 (.A(N586), .B(
        N594), .C(N601), .Y(ADD_32x32_fast_I271_un1_Y_0));
    NOR3A \off_div_RNIF00R1[14]  (.A(un1_off_divlto31_8), .B(
        off_div[16]), .C(off_div[14]), .Y(un1_off_divlto31_15));
    DFN1E0C0 \off_div[21]  (.D(\next_off_div[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[21]));
    XA1 \off_div_RNO[11]  (.A(N793), .B(ADD_32x32_fast_I301_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[11] ));
    XNOR2 un1_nsum_adj_I_40 (.A(sum_14), .B(N_11), .Y(I_40));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I42_Y (.A(off_div[24]), .B(
        off_div[25]), .C(sum_0_0), .Y(N488));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y (.A(
        ADD_32x32_fast_I263_un1_Y_0), .B(N796), .C(
        ADD_32x32_fast_I263_Y_1), .Y(N759));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I248_Y (.A(N654), .B(N538), 
        .C(N653), .Y(N799));
    NOR3A \off_div_RNIJNA01[30]  (.A(state[0]), .B(off_div[28]), .C(
        off_div[30]), .Y(next_off_div_2_sqmuxa_5));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I301_Y_0 (.A(sum_1_0), .B(
        \sum_adj[19]_net_1 ), .C(off_div[11]), .Y(
        ADD_32x32_fast_I301_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y (.A(
        ADD_32x32_fast_I260_un1_Y_0), .B(N787), .C(
        ADD_32x32_fast_I260_Y_2), .Y(N753));
    NOR2 \off_div_RNINVFT[12]  (.A(off_div[17]), .B(off_div[12]), .Y(
        un1_off_divlto31_8));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I306_Y_0 (.A(off_div[16]), 
        .B(sum_39), .Y(ADD_32x32_fast_I306_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I155_Y_0 (.A(off_div[29]), .B(
        off_div[30]), .C(sum_1_0), .Y(ADD_32x32_fast_I155_Y_0));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I80_Y (.A(N398), .B(
        off_div[6]), .C(\un1_sum_adj[6] ), .Y(N526));
    DFN1E1C0 \sum_adj[13]  (.D(\nsum_adj_5[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[13]_net_1 ));
    NOR3C \off_div_RNI6AFN5[14]  (.A(un1_off_divlto31_15), .B(
        un1_off_divlto31_14), .C(un1_off_divlto31_20), .Y(
        un1_off_divlto31_22));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I265_un1_Y_0 (.A(N624), .B(
        N640), .Y(ADD_32x32_fast_I265_un1_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I262_Y (.A(
        ADD_32x32_fast_I262_un1_Y_0), .B(N793), .C(
        ADD_32x32_fast_I262_Y_1), .Y(N757));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I170_Y (.A(N567), .B(N560), 
        .C(N559), .Y(N625));
    DFN1E0C0 \off_div[5]  (.D(\next_off_div[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[5]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I7_G0N (.A(\un1_sum_adj[7] )
        , .B(off_div[7]), .Y(N404));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I57_Y (.A(sum_1_0), .B(
        off_div[18]), .C(N435), .Y(N503));
    XOR2 \state_RNO[1]  (.A(state[1]), .B(state[0]), .Y(N_311_i));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I308_Y (.A(I236_un1_Y), .B(
        ADD_32x32_fast_I271_Y_0), .C(ADD_32x32_fast_I308_Y_0), .Y(
        \un1_off_div_1[18] ));
    MX2 \sum_adj_RNO[11]  (.A(sum_11), .B(I_32), .S(sum_1_0), .Y(
        \nsum_adj_5[11] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I321_Y_0 (.A(off_div[31]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I321_Y_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I116_Y (.A(N500), .B(N504), 
        .Y(N565));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I311_Y_0 (.A(off_div[21]), 
        .B(sum_39), .Y(ADD_32x32_fast_I311_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I269_Y_0 (.A(N647), .B(N632), 
        .C(N631), .Y(ADD_32x32_fast_I269_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I81_Y (.A(off_div[6]), .B(
        \un1_sum_adj[6] ), .C(N399), .Y(N527));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I245_Y (.A(N648), .B(N663), 
        .C(N647), .Y(N790));
    MX2 \sum_adj_RNO[12]  (.A(sum_12), .B(I_35), .S(sum_1_0), .Y(
        \nsum_adj_5[12] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I316_Y_0 (.A(off_div[26]), 
        .B(sum_39), .Y(ADD_32x32_fast_I316_Y_0));
    AND3 un1_nsum_adj_I_64 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[16] ), .Y(N_3));
    XOR2 \sum_adj_RNIC2OQ[17]  (.A(\sum_adj[17]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[9] ));
    AO1 \off_div_RNI732AB[31]  (.A(un1_off_divlto31_22), .B(
        un1_off_divlto31_21), .C(off_div[31]), .Y(next_off_div16));
    NOR3 un1_nsum_adj_I_67 (.A(sum_1_d0), .B(sum_0_d0), .C(sum_2_d0), 
        .Y(\DWACT_FINC_E[34] ));
    NOR2 \off_div_RNIT7IT[26]  (.A(off_div[27]), .B(off_div[26]), .Y(
        next_off_div_2_sqmuxa_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I70_Y (.A(N413), .B(N417), .C(
        N416), .Y(N516));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I192_Y (.A(N589), .B(N582), 
        .C(N581), .Y(N647));
    DFN1E0C0 \off_div[30]  (.D(\next_off_div[30] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[30]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I129_Y (.A(N513), .B(N517), 
        .Y(N578));
    XNOR2 un1_nsum_adj_I_46 (.A(sum_16), .B(N_9), .Y(I_46));
    NOR2A \state_RNIL6F5[0]  (.A(state[1]), .B(state[0]), .Y(
        \state_d[2] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I182_Y (.A(N579), .B(N572), 
        .C(N571), .Y(N637));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I127_Y (.A(N515), .B(N511), 
        .Y(N576));
    AND3 un1_nsum_adj_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_17));
    VCC VCC_i (.Y(VCC));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I249_Y (.A(I249_un1_Y), .B(
        N655), .Y(N802));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I0_G0N (.A(off_div[0]), .B(
        sum_2_0), .Y(N383));
    AND3 un1_nsum_adj_I_39 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[8] ), .Y(N_11));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I196_un1_Y (.A(N593), .B(
        N586), .Y(I196_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I45_Y (.A(off_div[23]), .B(
        off_div[24]), .C(sum_0_0), .Y(N491));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I111_Y (.A(N495), .B(N499), 
        .Y(N560));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I71_Y (.A(off_div[10]), .B(
        \un1_sum_adj[10] ), .C(N417), .Y(N517));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I9_G0N (.A(\un1_sum_adj[9] )
        , .B(off_div[9]), .Y(N410));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I228_un1_Y (.A(N643), .B(
        N628), .Y(I228_un1_Y));
    XOR2 \sum_adj_RNILF4N[20]  (.A(\sum_adj[20]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[12] ));
    NOR3B \state_RNIS9HFB_0[0]  (.A(state[1]), .B(state[0]), .C(
        next_off_div16), .Y(next_off_div_1_sqmuxa));
    XOR2 \sum_adj_RNISL3N[18]  (.A(\sum_adj[18]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[10] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I307_Y_0 (.A(off_div[17]), 
        .B(sum_39), .Y(ADD_32x32_fast_I307_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I2_G0N (.A(\un1_sum_adj[2] )
        , .B(off_div[2]), .Y(N389));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I148_Y (.A(N536), .B(N533), 
        .C(N532), .Y(N597));
    XOR2 \sum_adj_RNIB1OQ[16]  (.A(\sum_adj[16]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[8] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I48_Y (.A(off_div[22]), .B(
        off_div[21]), .C(sum_0_0), .Y(N494));
    NOR2 \off_div_RNIQ4IT[21]  (.A(off_div[21]), .B(off_div[29]), .Y(
        next_off_div_2_sqmuxa_4));
    NOR3C \off_div_RNIL71R1[17]  (.A(off_div[17]), .B(off_div[18]), .C(
        un5lto20_1), .Y(un5lto20_2));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I260_un1_Y_0 (.A(N614), .B(
        N630), .Y(ADD_32x32_fast_I260_un1_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I268_un1_Y (.A(N630), .B(
        N646), .C(N661), .Y(I268_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_3 (.A(N627), .B(N612), 
        .C(ADD_32x32_fast_I259_Y_2), .Y(ADD_32x32_fast_I259_Y_3));
    AO1C \state_RNIURLQM[1]  (.A(un5lt31), .B(next_off_div_2_sqmuxa_10)
        , .C(state[1]), .Y(un1_state_2_0));
    XNOR2 un1_nsum_adj_I_23 (.A(sum_8), .B(N_17), .Y(I_23_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I266_un1_Y_0 (.A(N642), .B(
        N626), .Y(ADD_32x32_fast_I266_un1_Y_0));
    XNOR2 un1_nsum_adj_I_28 (.A(sum_10), .B(N_15), .Y(I_28));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I67_Y (.A(off_div[13]), .B(
        \un1_sum_adj[13] ), .C(N420), .Y(N513));
    OR3 \off_div_RNI6NVQ1[11]  (.A(off_div[11]), .B(off_div[12]), .C(
        un5lto14_1), .Y(un5lto14_2));
    XNOR2 un1_nsum_adj_I_65 (.A(sum_22), .B(N_3), .Y(I_65));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I193_Y (.A(N590), .B(N582), 
        .Y(N648));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I5_G0N (.A(sum_1_0), .B(
        \sum_adj[13]_net_1 ), .C(off_div[5]), .Y(N398));
    AND3 un1_nsum_adj_I_52 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[12] ), .Y(N_7));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I317_Y_0 (.A(off_div[27]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I317_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y_1 (.A(N555), .B(N548), 
        .C(ADD_32x32_fast_I260_Y_0), .Y(ADD_32x32_fast_I260_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I243_Y (.A(N644), .B(N659), 
        .C(N643), .Y(N784));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I296_Y_0 (.A(off_div[6]), .B(
        \un1_sum_adj[6] ), .Y(ADD_32x32_fast_I296_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I183_Y (.A(N580), .B(N572), 
        .Y(N638));
    NOR3 un1_nsum_adj_I_60 (.A(sum_18), .B(sum_20), .C(sum_19), .Y(
        \DWACT_FINC_E[15] ));
    MX2 \sum_adj_RNO[8]  (.A(sum_8), .B(I_23_0), .S(sum_2_0), .Y(
        \nsum_adj_5[8] ));
    XA1 \off_div_RNO[6]  (.A(N659), .B(ADD_32x32_fast_I296_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[6] ));
    OR2 \off_div_RNILTFT[14]  (.A(off_div[13]), .B(off_div[14]), .Y(
        un5lto14_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I124_Y (.A(N512), .B(N509), 
        .C(N508), .Y(N573));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I273_Y_0 (.A(
        ADD_32x32_fast_I273_un1_Y_0), .B(N640), .C(N639), .Y(
        ADD_32x32_fast_I273_Y_0));
    NOR2 un1_nsum_adj_I_21 (.A(sum_6), .B(sum_7), .Y(\DWACT_FINC_E[3] )
        );
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I242_Y (.A(N642), .B(N657), 
        .C(N641), .Y(N781));
    DFN1E0C0 \off_div[1]  (.D(\next_off_div[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[1]));
    XA1 \off_div_RNO[8]  (.A(N802), .B(ADD_32x32_fast_I298_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[8] ));
    XNOR2 un1_nsum_adj_I_53 (.A(sum_18), .B(N_7), .Y(I_53));
    AND3 un1_nsum_adj_I_58 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[14] ), .Y(N_5));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I102_Y (.A(N490), .B(N486), 
        .Y(N551));
    OR2 \off_div_RNIJ4JA[3]  (.A(off_div[3]), .B(off_div[4]), .Y(
        un5lto4));
    MX2 \off_div_RNO[19]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[19] ), .S(\state_d_0[2] ), .Y(
        \next_off_div[19] ));
    DFN1E0C0 \off_div[10]  (.D(\next_off_div[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[10]));
    MX2 \off_div_RNO[10]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[10] ), .S(\state_d_0[2] ), .Y(
        \next_off_div[10] ));
    NOR3C \off_div_RNINOO35[6]  (.A(un1_off_divlto31_13), .B(
        un1_off_divlto31_12), .C(un1_off_divlto31_17), .Y(
        un1_off_divlto31_21));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I125_Y (.A(N509), .B(N513), 
        .Y(N574));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y_0 (.A(N553), .B(N561), 
        .Y(ADD_32x32_fast_I263_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I178_Y (.A(N575), .B(N568), 
        .C(N567), .Y(N633));
    DFN1E1C0 \sum_adj[12]  (.D(\nsum_adj_5[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[12]_net_1 ));
    XNOR2 un1_nsum_adj_I_49 (.A(sum_17), .B(N_8), .Y(I_49));
    MX2 \sum_adj_RNO[17]  (.A(sum_17), .B(I_49), .S(sum_2_0), .Y(
        \nsum_adj_5[17] ));
    NOR3A un1_nsum_adj_I_66 (.A(\DWACT_FINC_E[15] ), .B(sum_21), .C(
        sum_22), .Y(\DWACT_FINC_E[33] ));
    AND3 un1_nsum_adj_I_51 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[28] ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I297_Y (.A(\un1_sum_adj[7] ), 
        .B(off_div[7]), .C(N657), .Y(\un1_off_div_1[7] ));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I269_un1_Y (.A(N632), .B(
        N648), .C(N663), .Y(I269_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I136_Y (.A(N524), .B(N521), 
        .C(N520), .Y(N585));
    XA1 \off_div_RNO[16]  (.A(N779), .B(ADD_32x32_fast_I306_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[16] ));
    AO1C \state_RNIURLQM_0[1]  (.A(un5lt31), .B(
        next_off_div_2_sqmuxa_10), .C(state[1]), .Y(
        \state_RNIURLQM_0[1]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I35_Y (.A(off_div[29]), .B(
        off_div[28]), .C(sum_0_0), .Y(N481));
    MX2 \off_div_RNO[0]  (.A(next_off_div_0_sqmuxa), .B(
        \un1_off_div_1[0] ), .S(\state_d_0[2] ), .Y(\next_off_div[0] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I199_Y (.A(N596), .B(N588), 
        .Y(N654));
    XA1 \off_div_RNO[23]  (.A(N765), .B(ADD_32x32_fast_I313_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[23] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I264_un1_Y_0 (.A(N622), .B(
        N638), .Y(ADD_32x32_fast_I264_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I87_Y (.A(N393), .B(N390), 
        .Y(N533));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I189_Y (.A(N578), .B(N586), 
        .Y(N644));
    MX2 \off_div_RNO[18]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[18] ), .S(\state_d_0[2] ), .Y(
        \next_off_div[18] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I38_Y (.A(off_div[26]), .B(
        off_div[27]), .C(sum_0_0), .Y(N484));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I187_Y (.A(N576), .B(N584), 
        .Y(N642));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I273_Y (.A(N655), .B(N640), 
        .C(ADD_32x32_fast_I273_Y_0), .Y(N779));
    XA1 \off_div_RNO[25]  (.A(N761), .B(ADD_32x32_fast_I315_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[25] ));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I112_Y (.A(N500), .B(N496), 
        .Y(N561));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I14_G0N (.A(sum_0_0), .B(
        \sum_adj[22]_net_1 ), .C(off_div[14]), .Y(N425));
    DFN1E0C0 \off_div[12]  (.D(\next_off_div[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[12]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I271_Y_0 (.A(
        ADD_32x32_fast_I271_un1_Y_0), .B(N636), .C(N635), .Y(
        ADD_32x32_fast_I271_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I161_Y (.A(N485), .B(N489), 
        .C(N558), .Y(N616));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I103_Y (.A(N487), .B(N491), 
        .Y(N552));
    DFN1E0C0 \off_div[0]  (.D(\next_off_div[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[0]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I131_Y (.A(N515), .B(N519), 
        .Y(N580));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I120_Y (.A(N508), .B(N505), 
        .C(N504), .Y(N569));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I46_Y (.A(off_div[22]), .B(
        off_div[23]), .C(sum_0_0), .Y(N492));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I300_Y_0 (.A(off_div[10]), 
        .B(\un1_sum_adj[10] ), .Y(ADD_32x32_fast_I300_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I99_Y (.A(N483), .B(N487), 
        .Y(N548));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I77_Y (.A(off_div[8]), .B(
        \un1_sum_adj[8] ), .C(N405), .Y(N523));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I44_Y (.A(off_div[23]), .B(
        off_div[24]), .C(sum_0_0), .Y(N490));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y_2 (.A(N629), .B(N614), 
        .C(ADD_32x32_fast_I260_Y_1), .Y(ADD_32x32_fast_I260_Y_2));
    DFN1E1C0 \sum_adj[20]  (.D(\nsum_adj_5[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[20]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I53_Y (.A(off_div[20]), .B(
        off_div[19]), .C(sum_0_0), .Y(N499));
    MX2 \off_div_RNO[5]  (.A(next_off_div_0_sqmuxa), .B(
        \un1_off_div_1[5] ), .S(\state_d_0[2] ), .Y(\next_off_div[5] ));
    XA1 \off_div_RNO[2]  (.A(N601), .B(ADD_32x32_fast_I292_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[2] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I6_G0N (.A(\un1_sum_adj[6] )
        , .B(off_div[6]), .Y(N401));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I247_un1_Y (.A(N586), .B(
        N594), .C(N601), .Y(I247_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I151_Y (.A(N537), .B(
        \sum_adj_RNISG3M[8]_net_1 ), .C(N536), .Y(N601));
    XOR2 \sum_adj_RNIMG4N[21]  (.A(\sum_adj[21]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[13] ));
    DFN1E0P0 \off_div[6]  (.D(\next_off_div[6] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[6]));
    DFN1E1C0 \sum_adj[17]  (.D(\nsum_adj_5[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[17]_net_1 ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I320_Y_0 (.A(off_div[30]), 
        .B(sum_39), .Y(ADD_32x32_fast_I320_Y_0));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I305_Y (.A(\un1_sum_adj[15] )
        , .B(off_div[15]), .C(N781), .Y(\un1_off_div_1[15] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I310_Y_0 (.A(off_div[20]), 
        .B(sum_39), .Y(ADD_32x32_fast_I310_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I270_Y_0 (.A(N649), .B(N634), 
        .C(N633), .Y(ADD_32x32_fast_I270_Y_0));
    AND3 un1_nsum_adj_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E[4] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I230_un1_Y (.A(N645), .B(
        N630), .Y(I230_un1_Y));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I52_Y (.A(off_div[19]), .B(
        off_div[20]), .C(sum_0_0), .Y(N498));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I204_Y (.A(I204_un1_Y), .B(
        N595), .Y(N661));
    NOR3A un1_nsum_adj_I_27 (.A(\DWACT_FINC_E[4] ), .B(sum_8), .C(
        sum_9), .Y(N_15));
    NOR3A \off_div_RNID24R1[23]  (.A(un1_off_divlto31_4), .B(
        off_div[24]), .C(off_div[23]), .Y(un1_off_divlto31_13));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I263_un1_Y_0 (.A(N620), .B(
        N636), .Y(ADD_32x32_fast_I263_un1_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I194_Y (.A(N591), .B(N584), 
        .C(N583), .Y(N649));
    DFN1E0C0 \off_div[20]  (.D(\next_off_div[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[20]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I113_Y (.A(N501), .B(N497), 
        .Y(N562));
    OA1 \off_div_RNIGSN32[10]  (.A(un5lto9), .B(un5lt9), .C(
        off_div[10]), .Y(un5lt14));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I184_Y (.A(I184_un1_Y), .B(
        N573), .Y(N639));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_0 (.A(off_div[29]), .B(
        off_div[28]), .C(sum_1_0), .Y(ADD_32x32_fast_I259_Y_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I17_P0N (.A(off_div[17]), .B(
        sum_39), .Y(N435));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I294_Y_0 (.A(off_div[4]), .B(
        \un1_sum_adj[4] ), .Y(ADD_32x32_fast_I294_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I236_un1_Y (.A(N651), .B(
        N636), .Y(I236_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I10_G0N (.A(
        \un1_sum_adj[10] ), .B(off_div[10]), .Y(N413));
    XA1 \off_div_RNO[21]  (.A(N769), .B(ADD_32x32_fast_I311_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[21] ));
    DFN1E0C0 \off_div[18]  (.D(\next_off_div[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[18]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I262_un1_Y_0 (.A(N618), .B(
        N634), .Y(ADD_32x32_fast_I262_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I109_Y (.A(N493), .B(N497), 
        .Y(N558));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y_0 (.A(N486), .B(N482), 
        .Y(ADD_32x32_fast_I260_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I146_Y (.A(N534), .B(N531), 
        .C(N530), .Y(N595));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I107_Y (.A(N495), .B(N491), 
        .Y(N556));
    AND3 un1_nsum_adj_I_54 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[9] ), .C(\DWACT_FINC_E[12] ), .Y(
        \DWACT_FINC_E[13] ));
    AND3 un1_nsum_adj_I_69 (.A(\DWACT_FINC_E[29] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[33] ), .Y(N_2));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I195_Y (.A(N592), .B(N584), 
        .Y(N650));
    NOR2 un1_nsum_adj_I_57 (.A(sum_18), .B(sum_19), .Y(
        \DWACT_FINC_E[14] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I63_Y (.A(N429), .B(N426), 
        .Y(N509));
    NOR2A un1_nsum_adj_I_25 (.A(\DWACT_FINC_E[4] ), .B(sum_8), .Y(N_16)
        );
    NOR3A \off_div_RNINC4R1[27]  (.A(un1_off_divlto31_2), .B(
        off_div[27]), .C(off_div[28]), .Y(un1_off_divlto31_12));
    DFN1E0C0 \off_div[22]  (.D(\next_off_div[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[22]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I185_Y (.A(N574), .B(N582), 
        .Y(N640));
    NOR3C \off_div_RNI93FR2[24]  (.A(next_off_div_2_sqmuxa_2), .B(
        next_off_div_2_sqmuxa_1), .C(next_off_div_2_sqmuxa_5), .Y(
        next_off_div_2_sqmuxa_8));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I90_Y (.A(N383), .B(N387), .C(
        N386), .Y(N536));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I55_Y (.A(off_div[19]), .B(
        off_div[18]), .C(sum_0_0), .Y(N501));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I49_Y (.A(off_div[21]), .B(
        off_div[22]), .C(sum_0_0), .Y(N495));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_2 (.A(N553), .B(N546), 
        .C(ADD_32x32_fast_I259_Y_1), .Y(ADD_32x32_fast_I259_Y_2));
    XA1 \off_div_RNO[12]  (.A(N790), .B(ADD_32x32_fast_I302_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[12] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I62_Y (.A(N425), .B(N429), .C(
        N428), .Y(N508));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y (.A(
        ADD_32x32_fast_I261_un1_Y_0), .B(N790), .C(
        ADD_32x32_fast_I261_Y_2), .Y(N755));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I141_Y (.A(N529), .B(N525), 
        .Y(N590));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I36_Y (.A(off_div[28]), .B(
        off_div[27]), .C(sum_0_0), .Y(N482));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I7_P0N (.A(\un1_sum_adj[7] ), 
        .B(off_div[7]), .Y(N405));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I58_Y (.A(off_div[17]), .B(
        off_div[16]), .C(sum_1_0), .Y(N504));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I292_Y_0 (.A(off_div[2]), .B(
        \un1_sum_adj[2] ), .Y(ADD_32x32_fast_I292_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I91_Y (.A(sum_1_0), .B(
        off_div[0]), .C(N387), .Y(N537));
    DFN1E0C0 \off_div[17]  (.D(\next_off_div[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[17]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I119_Y (.A(N503), .B(N507), 
        .Y(N568));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I190_Y (.A(I190_un1_Y), .B(
        N579), .Y(N645));
    MX2 \sum_adj_RNO[23]  (.A(sum_23), .B(I_70), .S(sum_2_0), .Y(
        \nsum_adj_5[23] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I117_Y (.A(N501), .B(N505), 
        .Y(N566));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I132_Y (.A(N520), .B(N517), 
        .C(N516), .Y(N581));
    OA1 \off_div_RNI4T8N6[16]  (.A(off_div[16]), .B(un5lt16), .C(
        un5lto20_2), .Y(un5lt31));
    NOR3C \state_RNIS9HFB[0]  (.A(state[1]), .B(state[0]), .C(
        next_off_div16), .Y(next_off_div_0_sqmuxa));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I180_Y (.A(N577), .B(N570), 
        .C(N569), .Y(N635));
    NOR3B un1_nsum_adj_I_55 (.A(\DWACT_FINC_E[13] ), .B(
        \DWACT_FINC_E[28] ), .C(sum_18), .Y(N_6));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I128_Y (.A(N516), .B(N513), 
        .C(N512), .Y(N577));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I104_Y (.A(N492), .B(N488), 
        .Y(N553));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I9_P0N (.A(\un1_sum_adj[9] ), 
        .B(off_div[9]), .Y(N411));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I15_G0N (.A(
        \un1_sum_adj[15] ), .B(off_div[15]), .Y(N428));
    XOR2 \sum_adj_RNIOI4N[23]  (.A(\sum_adj[23]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[15] ));
    NOR3 un1_nsum_adj_I_50 (.A(sum_16), .B(sum_15), .C(sum_17), .Y(
        \DWACT_FINC_E[12] ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I295_Y_0 (.A(sum_1_0), .B(
        \sum_adj[13]_net_1 ), .C(off_div[5]), .Y(
        ADD_32x32_fast_I295_Y_0));
    XOR2 \sum_adj_RNI7TNQ[12]  (.A(\sum_adj[12]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[4] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I176_Y (.A(N573), .B(N566), 
        .C(N565), .Y(N631));
    XNOR2 un1_nsum_adj_I_26 (.A(sum_9), .B(N_16), .Y(I_26));
    NOR2 \off_div_RNIQ5JT[30]  (.A(off_div[30]), .B(off_div[29]), .Y(
        un1_off_divlto31_0));
    DFN1E0C0 \off_div[28]  (.D(\next_off_div[28] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[28]));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I83_Y (.A(off_div[4]), .B(
        \un1_sum_adj[4] ), .C(N399), .Y(N529));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I65_Y (.A(off_div[13]), .B(
        \un1_sum_adj[13] ), .C(N426), .Y(N511));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I12_P0N (.A(\un1_sum_adj[12] )
        , .B(off_div[12]), .Y(N420));
    DFN1C0 \state[1]  (.D(N_311_i), .CLK(clk_c), .CLR(n_rst_c), .Q(
        state[1]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I15_P0N (.A(\un1_sum_adj[15] )
        , .B(off_div[15]), .Y(N429));
    XA1 \off_div_RNO[31]  (.A(N749), .B(ADD_32x32_fast_I321_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[31] ));
    XA1 \off_div_RNO[14]  (.A(N784), .B(ADD_32x32_fast_I304_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[14] ));
    NOR2A \state_RNIL6F5_1[0]  (.A(state[0]), .B(state[1]), .Y(
        state_176_d));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I163_Y (.A(N552), .B(N560), 
        .Y(N618));
    NOR2 \off_div_RNIM0IT[21]  (.A(off_div[25]), .B(off_div[21]), .Y(
        un1_off_divlto31_4));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I133_Y (.A(N521), .B(N517), 
        .Y(N582));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I190_un1_Y (.A(N587), .B(
        N580), .Y(I190_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I68_Y (.A(N416), .B(N420), .C(
        N419), .Y(N514));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I114_Y (.A(N502), .B(N498), 
        .Y(N563));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I261_un1_Y_0 (.A(N616), .B(
        N632), .Y(ADD_32x32_fast_I261_un1_Y_0));
    XOR2 \sum_adj_RNIA0OQ[15]  (.A(\sum_adj[15]_net_1 ), .B(sum_2_0), 
        .Y(\un1_sum_adj[7] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I82_Y (.A(N395), .B(N399), .C(
        N398), .Y(N528));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I171_Y (.A(N560), .B(N568), 
        .Y(N626));
    NOR3 un1_nsum_adj_I_18 (.A(sum_3), .B(sum_5), .C(sum_4), .Y(
        \DWACT_FINC_E[2] ));
    MX2 \sum_adj_RNO[14]  (.A(sum_14), .B(I_40), .S(sum_2_0), .Y(
        \nsum_adj_5[14] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I40_Y (.A(off_div[25]), .B(
        off_div[26]), .C(sum_0_0), .Y(N486));
    DFN1E1C0 \sum_adj[8]  (.D(\nsum_adj_5[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[8]_net_1 ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I204_un1_Y (.A(N596), .B(
        N538), .Y(I204_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I12_G0N (.A(
        \un1_sum_adj[12] ), .B(off_div[12]), .Y(N419));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I11_P0N (.A(sum_1_0), .B(
        \sum_adj[19]_net_1 ), .C(off_div[11]), .Y(N417));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I73_Y (.A(off_div[10]), .B(
        \un1_sum_adj[10] ), .C(N411), .Y(N519));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I266_Y_0 (.A(N641), .B(N626), 
        .C(N625), .Y(ADD_32x32_fast_I266_Y_0));
    NOR3C \off_div_RNI44E12[5]  (.A(un1_off_divlto31_10), .B(
        un1_off_divlto31_9), .C(un1_off_divlt31), .Y(
        un1_off_divlto31_20));
    XNOR2 un1_nsum_adj_I_56 (.A(sum_19), .B(N_6), .Y(I_56));
    OA1B \state_RNO[0]  (.A(state[1]), .B(pwm_enable), .C(state[0]), 
        .Y(\state_ns[0] ));
    DFN1E0C0 \off_div[2]  (.D(\next_off_div[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[2]));
    NOR3C \off_div_RNIKUSF[5]  (.A(off_div[5]), .B(off_div[7]), .C(
        off_div[6]), .Y(un5lto7_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I39_Y (.A(off_div[27]), .B(
        off_div[26]), .C(sum_0_0), .Y(N485));
    DFN1E0C0 \off_div[27]  (.D(\next_off_div[27] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[27]));
    MX2 \sum_adj_RNO[18]  (.A(sum_18), .B(I_53), .S(sum_2_0), .Y(
        \nsum_adj_5[18] ));
    DFN1E1C0 \sum_adj[15]  (.D(\nsum_adj_5[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[15]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I41_Y (.A(off_div[26]), .B(
        off_div[25]), .C(sum_0_0), .Y(N487));
    XNOR2 un1_nsum_adj_I_32 (.A(sum_11), .B(N_14), .Y(I_32));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y (.A(
        ADD_32x32_fast_I264_un1_Y_0), .B(N799), .C(
        ADD_32x32_fast_I264_Y_1), .Y(N761));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I72_Y (.A(N410), .B(
        off_div[10]), .C(\un1_sum_adj[10] ), .Y(N518));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I295_Y (.A(
        ADD_32x32_fast_I295_Y_0), .B(N661), .Y(\un1_off_div_1[5] ));
    XA1 \off_div_RNO[29]  (.A(N753), .B(ADD_32x32_fast_I319_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[29] ));
    DFN1E0C0 \off_div[14]  (.D(\next_off_div[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[14]));
    DFN1E1C0 \sum_adj[10]  (.D(\nsum_adj_5[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[10]_net_1 ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I302_Y_0 (.A(off_div[12]), 
        .B(\un1_sum_adj[12] ), .Y(ADD_32x32_fast_I302_Y_0));
    MX2 \off_div_RNO[20]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[20] ), .S(\state_d_0[2] ), .Y(
        \next_off_div[20] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I300_Y (.A(
        ADD_32x32_fast_I300_Y_0), .B(N796), .Y(\un1_off_div_1[10] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I115_Y (.A(N503), .B(N499), 
        .Y(N564));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I258_un1_Y_0 (.A(N610), .B(
        N626), .Y(ADD_32x32_fast_I258_un1_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I142_Y (.A(N530), .B(N527), 
        .C(N526), .Y(N591));
    NOR2 \off_div_RNIHPFT[10]  (.A(off_div[13]), .B(off_div[10]), .Y(
        un1_off_divlto31_9));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I56_Y (.A(off_div[17]), .B(
        off_div[18]), .C(sum_0_0), .Y(N502));
    XA1 \off_div_RNO[26]  (.A(N759), .B(ADD_32x32_fast_I316_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[26] ));
    MX2 \sum_adj_RNO[13]  (.A(sum_13), .B(I_37), .S(sum_1_0), .Y(
        \nsum_adj_5[13] ));
    DFN1E1C0 \sum_adj[19]  (.D(\nsum_adj_5[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[19]_net_1 ));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I267_un1_Y (.A(N628), .B(
        N644), .C(N659), .Y(I267_un1_Y));
    MX2 \off_div_RNO[17]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[17] ), .S(\state_d_0[2] ), .Y(
        \next_off_div[17] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I54_Y (.A(off_div[18]), .B(
        off_div[19]), .C(sum_0_0), .Y(N500));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I267_Y (.A(I228_un1_Y), .B(
        N627), .C(I267_un1_Y), .Y(N767));
    NOR2 \off_div_RNIS4GT[15]  (.A(off_div[19]), .B(off_div[15]), .Y(
        un1_off_divlto31_6));
    DFN1E0C0 \off_div[4]  (.D(\next_off_div[4] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[4]));
    NOR3 un1_nsum_adj_I_33 (.A(sum_10), .B(sum_9), .C(sum_11), .Y(
        \DWACT_FINC_E[7] ));
    NOR2 un1_nsum_adj_I_38 (.A(sum_12), .B(sum_13), .Y(
        \DWACT_FINC_E[8] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I303_Y_0 (.A(off_div[13]), 
        .B(\un1_sum_adj[13] ), .Y(ADD_32x32_fast_I303_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I169_Y (.A(N558), .B(N566), 
        .Y(N624));
    DFN1E0C0 \off_div[19]  (.D(\next_off_div[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[19]));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I85_Y (.A(off_div[4]), .B(
        \un1_sum_adj[4] ), .C(N393), .Y(N531));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I312_Y_0 (.A(off_div[22]), 
        .B(sum_39), .Y(ADD_32x32_fast_I312_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I139_Y (.A(N527), .B(N523), 
        .Y(N588));
    XA1 \off_div_RNO[28]  (.A(N755), .B(ADD_32x32_fast_I318_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[28] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I167_Y (.A(N564), .B(N556), 
        .Y(N622));
    DFN1E0C0 \off_div[16]  (.D(\next_off_div[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[16]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I198_Y (.A(N595), .B(N588), 
        .C(N587), .Y(N653));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I137_Y (.A(N521), .B(N525), 
        .Y(N586));
    DFN1E0C0 \off_div[8]  (.D(\next_off_div[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[8]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I97_Y (.A(N485), .B(N481), 
        .Y(N546));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I188_Y (.A(N585), .B(N578), 
        .C(N577), .Y(N643));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I16_P0N (.A(off_div[16]), .B(
        sum_39), .Y(N432));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I110_Y (.A(N494), .B(N498), 
        .Y(N559));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I88_Y (.A(N386), .B(N390), .C(
        N389), .Y(N534));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0 (.A(off_div[30]), .B(
        off_div[29]), .C(sum_1_0), .Y(ADD_32x32_fast_I258_Y_0));
    NOR3 un1_nsum_adj_I_29 (.A(sum_7), .B(sum_6), .C(sum_8), .Y(
        \DWACT_FINC_E[5] ));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I310_Y (.A(I269_un1_Y), .B(
        ADD_32x32_fast_I269_Y_0), .C(ADD_32x32_fast_I310_Y_0), .Y(
        \un1_off_div_1[20] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y_2 (.A(N616), .B(N631), 
        .C(ADD_32x32_fast_I261_Y_1), .Y(ADD_32x32_fast_I261_Y_2));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I159_Y (.A(N556), .B(N548), 
        .Y(N614));
    NOR3A un1_nsum_adj_I_31 (.A(\DWACT_FINC_E[6] ), .B(sum_9), .C(
        sum_10), .Y(N_14));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I313_Y_0 (.A(off_div[23]), 
        .B(sum_39), .Y(ADD_32x32_fast_I313_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I157_Y (.A(N489), .B(N493), 
        .C(N546), .Y(N612));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I75_Y (.A(off_div[8]), .B(
        \un1_sum_adj[8] ), .C(N411), .Y(N521));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I293_Y (.A(
        ADD_32x32_fast_I293_Y_0), .B(N599), .Y(\un1_off_div_1[3] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I143_Y (.A(N531), .B(N527), 
        .Y(N592));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I259_un1_Y_0 (.A(N612), .B(
        N628), .Y(ADD_32x32_fast_I259_un1_Y_0));
    DFN1E0P0 \off_div[3]  (.D(\next_off_div[3] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[3]));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I290_Y (.A(sum_2_0), .B(
        off_div[0]), .C(\sum_adj_RNISG3M[8]_net_1 ), .Y(
        \un1_off_div_1[0] ));
    MX2 \off_div_RNO[7]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[7] ), .S(\state_d_0[2] ), .Y(\next_off_div[7] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I78_Y (.A(N401), .B(N405), .C(
        N404), .Y(N524));
    DFN1E1C0 \sum_adj[21]  (.D(\nsum_adj_5[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[21]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_3 (.A(N610), .B(N625), 
        .C(ADD_32x32_fast_I258_Y_2), .Y(ADD_32x32_fast_I258_Y_3));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I66_Y (.A(N419), .B(
        off_div[13]), .C(\un1_sum_adj[13] ), .Y(N512));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I270_un1_Y (.A(N634), .B(
        N650), .C(N599), .Y(I270_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I8_G0N (.A(\un1_sum_adj[8] )
        , .B(off_div[8]), .Y(N407));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I224_un1_Y (.A(N639), .B(
        N624), .Y(I224_un1_Y));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I299_Y_0 (.A(off_div[9]), .B(
        \un1_sum_adj[9] ), .Y(ADD_32x32_fast_I299_Y_0));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I1_G0N (.A(sum_1_0), .B(
        \sum_adj[9]_net_1 ), .C(off_div[1]), .Y(N386));
    XA1 \off_div_RNO[4]  (.A(N663), .B(ADD_32x32_fast_I294_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[4] ));
    DFN1E0C0 \off_div[24]  (.D(\next_off_div[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNIURLQM_0[1]_net_1 ), .Q(off_div[24]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I64_Y (.A(N422), .B(N426), .C(
        N425), .Y(N510));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I205_Y (.A(N598), .B(
        \sum_adj_RNISG3M[8]_net_1 ), .C(N597), .Y(N663));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I172_Y (.A(N569), .B(N562), 
        .C(N561), .Y(N627));
    XNOR2 un1_nsum_adj_I_59 (.A(sum_20), .B(N_5), .Y(I_59));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I3_G0N (.A(sum_1_0), .B(
        \sum_adj[11]_net_1 ), .C(off_div[3]), .Y(N392));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I134_Y (.A(N522), .B(N519), 
        .C(N518), .Y(N583));
    AND3 un1_nsum_adj_I_42 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[9] ), .Y(N_10));
    DFN1E1C0 \sum_adj[16]  (.D(\nsum_adj_5[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[16]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I244_Y (.A(N646), .B(N661), 
        .C(N645), .Y(N787));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I238_un1_Y (.A(N653), .B(
        N638), .Y(I238_un1_Y));
    MX2 \sum_adj_RNO[19]  (.A(sum_19), .B(I_56), .S(sum_2_0), .Y(
        \nsum_adj_5[19] ));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y_1 (.A(N488), .B(N484), 
        .C(N557), .Y(ADD_32x32_fast_I261_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I126_Y (.A(N514), .B(N511), 
        .C(N510), .Y(N575));
    NOR2A \state_RNIL6F5_0[0]  (.A(state[1]), .B(state[0]), .Y(
        \state_d_0[2] ));
    XA1 \off_div_RNO[30]  (.A(N751), .B(ADD_32x32_fast_I320_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[30] ));
    
endmodule


module integral_calc_13s_4(
       avg_old,
       avg_new,
       LED_33,
       LED_FB,
       LED_5,
       LED_c,
       LED_15,
       choose,
       choose_0_0,
       LED_12,
       average,
       LED_12_i_0,
       avg_done,
       calc_avg,
       n_rst_c,
       clk_c
    );
input  [11:0] avg_old;
input  [11:0] avg_new;
input  [7:6] LED_33;
input  [7:6] LED_FB;
input  [7:6] LED_5;
output [7:6] LED_c;
input  [7:6] LED_15;
input  [2:0] choose;
input  choose_0_0;
output [7:0] LED_12;
output [6:2] average;
output LED_12_i_0;
output avg_done;
input  calc_avg;
input  n_rst_c;
input  clk_c;

    wire \state_1[0]_net_1 , \state_1_RNI4F701[0]_net_1 , 
        \state_0[0]_net_1 , avg_done_0, \state[1]_net_1 , 
        ADD_26x26_fast_I253_Y_0, \integ[23]_net_1 , \state[0]_net_1 , 
        ADD_26x26_fast_I254_Y_0, \integ[24]_net_1 , 
        ADD_26x26_fast_I255_Y_0, \integ[25]_net_1 , 
        ADD_26x26_fast_I206_Y_2, N506, N521, ADD_26x26_fast_I206_Y_1, 
        N452, N459, ADD_26x26_fast_I206_Y_0, N402, N398, 
        ADD_26x26_fast_I252_Y_0, \integ[22]_net_1 , 
        ADD_26x26_fast_I204_Y_3, N502, N517, ADD_26x26_fast_I204_Y_2, 
        ADD_26x26_fast_I204_Y_0, N455, ADD_26x26_fast_I205_Y_3, N504, 
        N519, ADD_26x26_fast_I205_Y_2, N400, ADD_26x26_fast_I205_Y_0, 
        N457, ADD_26x26_fast_I251_Y_0, \integ[21]_net_1 , 
        ADD_26x26_fast_I250_Y_0, \integ[20]_net_1 , 
        ADD_26x26_fast_I249_Y_0, \integ[19]_net_1 , 
        ADD_26x26_fast_I207_Y_2, N508, N523, ADD_26x26_fast_I207_Y_1, 
        N461, N454, ADD_26x26_fast_I207_Y_0, N404, 
        ADD_26x26_fast_I206_un1_Y_0, N522, ADD_26x26_fast_I246_Y_0, 
        \integ[16]_net_1 , ADD_26x26_fast_I247_Y_0, \integ[17]_net_1 , 
        ADD_26x26_fast_I248_Y_0, \integ[18]_net_1 , 
        ADD_26x26_fast_I241_Y_0, \un18_next_int_m[11] , 
        \inf_abs0_m[11] , ADD_26x26_fast_I208_Y_1, 
        ADD_26x26_fast_I208_un1_Y_0, N541, ADD_26x26_fast_I208_Y_0, 
        N463, N456, ADD_26x26_fast_I209_Y_1, 
        ADD_26x26_fast_I209_un1_Y_0, N543, ADD_26x26_fast_I209_Y_0, 
        N465, N458, ADD_26x26_fast_I239_Y_0, \un18_next_int_m[9] , 
        \inf_abs0_m[9] , ADD_26x26_fast_I238_Y_0, \un1_next_int[8] , 
        ADD_26x26_fast_I210_Y_1, ADD_26x26_fast_I210_un1_Y_0, N491, 
        ADD_26x26_fast_I210_Y_0, N467, N460, 
        ADD_26x26_fast_I205_un1_Y_0, N520, ADD_26x26_fast_I204_un1_Y_0, 
        N518, ADD_26x26_fast_I240_Y_0, \state_1_RNIH8S81[0]_net_1 , 
        ADD_26x26_fast_I212_Y_0, ADD_26x26_fast_I212_un1_Y_0, 
        ADD_26x26_fast_I211_Y_1, ADD_26x26_fast_I211_un1_Y_0, N532, 
        ADD_26x26_fast_I211_Y_0, N469, N462, ADD_26x26_fast_I213_Y_0, 
        ADD_26x26_fast_I213_un1_Y_0, ADD_26x26_fast_I234_Y_0, 
        \state_RNI72LK1[0]_net_1 , ADD_26x26_fast_I235_Y_0, 
        \inf_abs0_m[5] , \un18_next_int_m[5] , N512, N528, N510, N526, 
        N476, N484, N514, N488, N480, N442, N482, N490, 
        \state_1_RNIF5VI1[0]_net_1 , N470, N493, 
        ADD_26x26_fast_I232_Y_0, \state_RNI3UKK1[0]_net_1 , 
        ADD_26x26_fast_I231_Y_0, \un18_next_int_m[1] , \inf_abs0_m[1] , 
        \integ[1]_net_1 , ADD_26x26_fast_I127_Y_0, 
        ADD_26x26_fast_I125_Y_0, ADD_26x26_fast_I230_Y_0, 
        \integ[0]_net_1 , \un1_integ[21] , I176_un1_Y, \un1_integ[17] , 
        I184_un1_Y, \un1_integ[12] , N646, I207_un1_Y, N524, N539, 
        \un1_integ[20] , I178_un1_Y, \un1_integ[22] , \un1_integ[19] , 
        I180_un1_Y, \un1_integ[3] , \state_RNI50LK1[0]_net_1 , 
        \un1_integ[18] , I182_un1_Y, \un1_integ[25] , I204_un1_Y, 
        \un1_integ[6] , \state_RNIB6LK1[0]_net_1 , \un1_integ[14] , 
        N640, \un1_integ[16] , I186_un1_Y, \un1_integ[24] , I205_un1_Y, 
        \un1_integ[0] , \un1_integ[7] , \state_RNID8LK1[0]_net_1 , 
        N537, \un1_integ[13] , N643, \un1_integ[15] , 
        \integ[15]_net_1 , N637, \un1_integ[23] , I206_un1_Y, 
        \un1_integ[2] , \un1_integ[10] , N531, I193_un1_Y, 
        \un1_integ[11] , N529, I192_un1_Y, \un1_integ[9] , N533, 
        I194_un1_Y, \un1_integ[8] , N535, I195_un1_Y, \un1_integ[5] , 
        \un1_integ[4] , \un1_integ[1] , N401, N399, N474, N489, N481, 
        I163_un1_Y, N439, N435, N330, N321, N324, N527, N473, N477, 
        N466, N464, N411, N415, N471, N440, N437, N436, N323, N441, 
        N318, N429, N433, N333, I74_un1_Y, N317, N468, N419, N422, 
        N418, N483, N431, N434, N430, N487, N438, N475, I148_un1_Y, 
        N479, N472, N525, I152_un1_Y, I160_un1_Y, N486, N414, N320, 
        N326, N329, I121_un1_Y, N485, N478, N342, N341, N407, 
        I162_un1_Y, N408, N410, N405, N_65, N_57, N_41, N_49, N_73, 
        N_104, N403, N406, \inf_abs0_m[8] , \un18_next_int_m[8] , 
        N_103, N_48, N_40, N_72, N_56, N_64, N426, N338, N427, N424, 
        N421, N420, N347, N351, N350, N348, N425, N345, N417, N416, 
        N336, N413, N423, N428, N335, N344, \inf_abs0_m[0] , 
        \un18_next_int_m[0] , \inf_abs0_m[3] , \un18_next_int_m[3] , 
        \inf_abs0_m[4] , \un18_next_int_m[4] , \inf_abs0_m[7] , 
        \un18_next_int_m[7] , \inf_abs0_m[10] , \un18_next_int_m[10] , 
        \inf_abs0_m[2] , \un18_next_int_m[2] , \inf_abs0_m[6] , 
        \un18_next_int_m[6] , \state_RNO[1]_net_1 , N412, N409, N354, 
        N353, N357, N332, N432, GND, VCC;
    
    AO1 un1_integ_0_0_ADD_26x26_fast_I56_Y (.A(N341), .B(N345), .C(
        N344), .Y(N424));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I148_un1_Y (.A(N479), .B(N472), 
        .Y(I148_un1_Y));
    NOR2 \state_0_RNIO46P[0]  (.A(\state[1]_net_1 ), .B(
        \state_0[0]_net_1 ), .Y(avg_done_0));
    MX2 \un1_integ_0_0_LED_7[7]  (.A(N_49), .B(N_73), .S(choose[0]), 
        .Y(LED_c[7]));
    DFN1C0 \state[0]  (.D(\state_1_RNI4F701[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state[0]_net_1 ));
    DFN1E0C0 \integ[13]  (.D(\un1_integ[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_12[6]));
    DFN1E0C0 \integ[24]  (.D(\un1_integ[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[24]_net_1 ));
    NOR2A \state_RNIKNMQ[1]  (.A(\state[1]_net_1 ), .B(avg_old[2]), .Y(
        \un18_next_int_m[2] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I61_Y (.A(
        \state_RNID8LK1[0]_net_1 ), .B(LED_12[0]), .C(N336), .Y(N429));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I248_Y_0 (.A(\integ[18]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I248_Y_0));
    NOR2A \state_RNIILMQ[1]  (.A(\state[1]_net_1 ), .B(avg_old[0]), .Y(
        \un18_next_int_m[0] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I41_Y (.A(\integ[17]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N409));
    NOR2A \state_RNIRUMQ[1]  (.A(\state[1]_net_1 ), .B(avg_old[9]), .Y(
        \un18_next_int_m[9] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I204_un1_Y (.A(N533), .B(
        I194_un1_Y), .C(ADD_26x26_fast_I204_un1_Y_0), .Y(I204_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I86_Y (.A(N404), .B(N408), .Y(
        N457));
    NOR2B \state_RNIF6UP[0]  (.A(avg_new[2]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[2] ));
    MX2 \un1_integ_0_0_LED_7[6]  (.A(N_48), .B(N_72), .S(choose[0]), 
        .Y(LED_c[6]));
    NOR2B \state_RNIJAUP[0]  (.A(avg_new[6]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[6] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I98_Y (.A(N420), .B(N417), .C(
        N416), .Y(N469));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I176_un1_Y (.A(N510), .B(N525), 
        .Y(I176_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I205_un1_Y_0 (.A(N504), .B(N520)
        , .Y(ADD_26x26_fast_I205_un1_Y_0));
    NOR2A \un1_integ_0_0_LED_5[6]  (.A(LED_33[6]), .B(choose[2]), .Y(
        N_64));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I51_Y (.A(N354), .B(N351), .Y(
        N419));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y (.A(
        ADD_26x26_fast_I230_Y_0), .B(\state_1_RNIF5VI1[0]_net_1 ), .Y(
        \un1_integ[0] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I253_Y (.A(I206_un1_Y), .B(
        ADD_26x26_fast_I206_Y_2), .C(ADD_26x26_fast_I253_Y_0), .Y(
        \un1_integ[23] ));
    DFN1E0C0 \integ[21]  (.D(\un1_integ[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[21]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I146_Y (.A(N470), .B(N477), .C(
        N469), .Y(N523));
    NOR2B \state_1_RNIUG8O[0]  (.A(avg_new[1]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[1] ));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I210_un1_Y_0 (.A(N476), .B(N484)
        , .C(N514), .Y(ADD_26x26_fast_I210_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I142_Y (.A(N473), .B(N466), .C(
        N465), .Y(N519));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I231_Y (.A(
        ADD_26x26_fast_I231_Y_0), .B(N442), .Y(\un1_integ[1] ));
    NOR2B \state_RNII9UP[0]  (.A(avg_new[5]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[5] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I155_Y (.A(N486), .B(N478), .Y(
        N532));
    DFN1E0C0 \integ[15]  (.D(\un1_integ[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[15]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I103_Y (.A(N425), .B(N421), .Y(
        N474));
    NOR2B \state_1_RNIEVUM[0]  (.A(avg_new[10]), .B(\state_1[0]_net_1 )
        , .Y(\inf_abs0_m[10] ));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I125_Y (.A(N399), .B(
        ADD_26x26_fast_I125_Y_0), .C(N456), .Y(N502));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_1 (.A(
        ADD_26x26_fast_I209_un1_Y_0), .B(N543), .C(
        ADD_26x26_fast_I209_Y_0), .Y(ADD_26x26_fast_I209_Y_1));
    MX2 \un1_integ_0_0_LED_1[6]  (.A(LED_12[6]), .B(LED_15[6]), .S(
        choose_0_0), .Y(N_103));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I97_Y (.A(N419), .B(N415), .Y(
        N468));
    AO1 un1_integ_0_0_ADD_26x26_fast_I94_Y (.A(N416), .B(N413), .C(
        N412), .Y(N465));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I81_Y (.A(N403), .B(N399), .Y(
        N452));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I151_Y (.A(N474), .B(N482), .Y(
        N528));
    OR2 un1_integ_0_0_ADD_26x26_fast_I74_Y (.A(I74_un1_Y), .B(N317), 
        .Y(N442));
    AX1D un1_integ_0_0_ADD_26x26_fast_I238_Y (.A(N535), .B(I195_un1_Y), 
        .C(ADD_26x26_fast_I238_Y_0), .Y(\un1_integ[8] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I121_Y (.A(I121_un1_Y), .B(N440), 
        .Y(N493));
    AO1 un1_integ_0_0_ADD_26x26_fast_I190_Y (.A(N526), .B(N541), .C(
        N525), .Y(N643));
    NOR2A \state_RNINQMQ[1]  (.A(\state[1]_net_1 ), .B(avg_old[5]), .Y(
        \un18_next_int_m[5] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I5_P0N (.A(\inf_abs0_m[5] ), .B(
        \un18_next_int_m[5] ), .C(average[5]), .Y(N333));
    NOR2A \state_RNIORMQ[1]  (.A(\state[1]_net_1 ), .B(avg_old[6]), .Y(
        \un18_next_int_m[6] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I246_Y (.A(I186_un1_Y), .B(
        ADD_26x26_fast_I213_Y_0), .C(ADD_26x26_fast_I246_Y_0), .Y(
        \un1_integ[16] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I252_Y_0 (.A(\integ[22]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I252_Y_0));
    DFN1C0 \state_1[0]  (.D(\state_1_RNI4F701[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_1[0]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I39_Y (.A(\integ[18]_net_1 ), .B(
        \integ[17]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N407));
    OA1B un1_integ_0_0_ADD_26x26_fast_I32_Y (.A(\integ[20]_net_1 ), .B(
        \integ[21]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N400));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I194_un1_Y (.A(N488), .B(N480), 
        .C(N442), .Y(I194_un1_Y));
    AO1B un1_integ_0_0_ADD_26x26_fast_I125_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\integ[24]_net_1 ), .C(\state_1[0]_net_1 ), .Y(
        ADD_26x26_fast_I125_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I100_Y (.A(N422), .B(N419), .C(
        N418), .Y(N471));
    OR2 un1_integ_0_0_ADD_26x26_fast_I12_P0N (.A(LED_12[5]), .B(
        \state[1]_net_1 ), .Y(N354));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I10_G0N (.A(LED_12[3]), .B(
        \state_1_RNIH8S81[0]_net_1 ), .Y(N347));
    DFN1E0C0 \integ[12]  (.D(\un1_integ[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_12[5]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I109_Y (.A(N431), .B(N427), .Y(
        N480));
    OA1B un1_integ_0_0_ADD_26x26_fast_I205_Y_0 (.A(\integ[22]_net_1 ), 
        .B(\integ[23]_net_1 ), .C(\state_1[0]_net_1 ), .Y(
        ADD_26x26_fast_I205_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I115_Y (.A(N433), .B(N437), .Y(
        N486));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I12_G0N (.A(LED_12[5]), .B(
        \state[1]_net_1 ), .Y(N353));
    MX2 \un1_integ_0_0_LED_3[6]  (.A(N_103), .B(N_40), .S(choose[1]), 
        .Y(N_48));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_0 (.A(N463), .B(N456), .C(
        N455), .Y(ADD_26x26_fast_I208_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I111_Y (.A(N429), .B(N433), .Y(
        N482));
    OR2 un1_integ_0_0_ADD_26x26_fast_I2_P0N (.A(
        \state_RNI3UKK1[0]_net_1 ), .B(average[2]), .Y(N324));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I250_Y_0 (.A(\integ[20]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I250_Y_0));
    DFN1E0C0 \integ[10]  (.D(\un1_integ[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_12[3]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I180_un1_Y (.A(N514), .B(N529), 
        .Y(I180_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I162_Y (.A(I162_un1_Y), .B(N487), 
        .Y(N541));
    NOR2A \un1_integ_0_0_LED_2[6]  (.A(LED_5[6]), .B(choose_0_0), .Y(
        N_40));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I6_G0N (.A(average[6]), .B(
        \state_RNIB6LK1[0]_net_1 ), .Y(N335));
    INV \integ_RNITE71[12]  (.A(LED_12[5]), .Y(LED_12_i_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I249_Y (.A(I180_un1_Y), .B(
        ADD_26x26_fast_I210_Y_1), .C(ADD_26x26_fast_I249_Y_0), .Y(
        \un1_integ[19] ));
    GND GND_i (.Y(GND));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I246_Y_0 (.A(\integ[16]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I246_Y_0));
    NOR2B \state_RNIMDUP[0]  (.A(avg_new[9]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[9] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I6_P0N (.A(average[6]), .B(
        \state_RNIB6LK1[0]_net_1 ), .Y(N336));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I212_un1_Y_0 (.A(N488), .B(N480)
        , .C(N442), .Y(ADD_26x26_fast_I212_un1_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I1_G0N (.A(\un18_next_int_m[1] ), 
        .B(\inf_abs0_m[1] ), .C(\integ[1]_net_1 ), .Y(N320));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I107_Y (.A(N429), .B(N425), .Y(
        N478));
    OA1B un1_integ_0_0_ADD_26x26_fast_I38_Y (.A(\integ[17]_net_1 ), .B(
        \integ[18]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N406));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I209_un1_Y_0 (.A(N512), .B(N528)
        , .Y(ADD_26x26_fast_I209_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_3 (.A(N504), .B(N519), .C(
        ADD_26x26_fast_I205_Y_2), .Y(ADD_26x26_fast_I205_Y_3));
    AX1D un1_integ_0_0_ADD_26x26_fast_I255_Y (.A(I204_un1_Y), .B(
        ADD_26x26_fast_I204_Y_3), .C(ADD_26x26_fast_I255_Y_0), .Y(
        \un1_integ[25] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I204_Y_0 (.A(\integ[24]_net_1 ), 
        .B(\integ[23]_net_1 ), .C(\state_1[0]_net_1 ), .Y(
        ADD_26x26_fast_I204_Y_0));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I243_Y (.A(\state_1[0]_net_1 ), 
        .B(LED_12[6]), .C(N643), .Y(\un1_integ[13] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I231_Y_0 (.A(
        \un18_next_int_m[1] ), .B(\inf_abs0_m[1] ), .C(
        \integ[1]_net_1 ), .Y(ADD_26x26_fast_I231_Y_0));
    NOR2A \state_RNIJMMQ[1]  (.A(\state[1]_net_1 ), .B(avg_old[1]), .Y(
        \un18_next_int_m[1] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I69_Y (.A(average[3]), .B(
        \state_RNI50LK1[0]_net_1 ), .C(N324), .Y(N437));
    AO1 un1_integ_0_0_ADD_26x26_fast_I62_Y (.A(N332), .B(N336), .C(
        N335), .Y(N430));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I193_un1_Y (.A(N532), .B(N493), 
        .Y(I193_un1_Y));
    NOR2B \state_RNILCUP[0]  (.A(avg_new[8]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[8] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I152_un1_Y (.A(N483), .B(N476), 
        .Y(I152_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I7_G0N (.A(LED_12[0]), .B(
        \state_RNID8LK1[0]_net_1 ), .Y(N338));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I49_Y (.A(N357), .B(N354), .Y(
        N417));
    OA1B un1_integ_0_0_ADD_26x26_fast_I42_Y (.A(\integ[15]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N410));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I145_Y (.A(N476), .B(N468), .Y(
        N522));
    OR2 un1_integ_0_0_ADD_26x26_fast_I10_P0N (.A(LED_12[3]), .B(
        \state_1_RNIH8S81[0]_net_1 ), .Y(N348));
    OR3 un1_integ_0_0_ADD_26x26_fast_I1_P0N (.A(\un18_next_int_m[1] ), 
        .B(\inf_abs0_m[1] ), .C(\integ[1]_net_1 ), .Y(N321));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I184_un1_Y (.A(N533), .B(N518), 
        .Y(I184_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I192_un1_Y (.A(N476), .B(N484), 
        .C(N491), .Y(I192_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I141_Y (.A(N464), .B(N472), .Y(
        N518));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I93_Y (.A(N411), .B(N415), .Y(
        N464));
    AO1B un1_integ_0_0_ADD_26x26_fast_I37_Y (.A(\integ[18]_net_1 ), .B(
        \integ[19]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N405));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I0_G0N (.A(\integ[0]_net_1 ), 
        .B(\state[1]_net_1 ), .Y(N317));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I73_Y (.A(N318), .B(N321), .Y(
        N441));
    OA1 un1_integ_0_0_ADD_26x26_fast_I59_Y (.A(
        \state_RNID8LK1[0]_net_1 ), .B(LED_12[0]), .C(N342), .Y(N427));
    AO1 un1_integ_0_0_ADD_26x26_fast_I52_Y (.A(N347), .B(N351), .C(
        N350), .Y(N420));
    NOR2A \state_RNO[1]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 ), 
        .Y(\state_RNO[1]_net_1 ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I34_Y (.A(\integ[19]_net_1 ), .B(
        \integ[20]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N402));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I236_Y (.A(
        \state_RNIB6LK1[0]_net_1 ), .B(average[6]), .C(N539), .Y(
        \un1_integ[6] ));
    OR2 \state_1_RNIH8S81[0]  (.A(\inf_abs0_m[10] ), .B(
        \un18_next_int_m[10] ), .Y(\state_1_RNIH8S81[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I150_Y (.A(N481), .B(N474), .C(
        N473), .Y(N527));
    DFN1E0C0 \integ[0]  (.D(\un1_integ[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(\integ[0]_net_1 ));
    NOR3A \state_1_RNI4F701[0]  (.A(calc_avg), .B(\state[1]_net_1 ), 
        .C(\state_1[0]_net_1 ), .Y(\state_1_RNI4F701[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I120_Y (.A(N439), .B(N442), .C(
        N438), .Y(N491));
    AO1 un1_integ_0_0_ADD_26x26_fast_I104_Y (.A(N426), .B(N423), .C(
        N422), .Y(N475));
    NOR2B \state_RNIG7UP[0]  (.A(avg_new[3]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[3] ));
    VCC VCC_i (.Y(VCC));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I129_Y (.A(N452), .B(N460), .Y(
        N506));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I113_Y (.A(N431), .B(N435), .Y(
        N484));
    AX1D un1_integ_0_0_ADD_26x26_fast_I241_Y_0 (.A(
        \un18_next_int_m[11] ), .B(\inf_abs0_m[11] ), .C(LED_12[4]), 
        .Y(ADD_26x26_fast_I241_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I89_Y (.A(N407), .B(N411), .Y(
        N460));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I68_Y (.A(N323), .B(average[3]), 
        .C(\state_RNI50LK1[0]_net_1 ), .Y(N436));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_0 (.A(N469), .B(N462), .C(
        N461), .Y(ADD_26x26_fast_I211_Y_0));
    NOR2A \un1_integ_0_0_LED_4[7]  (.A(LED_FB[7]), .B(choose[2]), .Y(
        N_57));
    DFN1E0C0 \integ[4]  (.D(\un1_integ[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[4]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I108_Y (.A(N430), .B(N427), .C(
        N426), .Y(N479));
    NOR2A \state_RNIMPMQ[1]  (.A(\state[1]_net_1 ), .B(avg_old[4]), .Y(
        \un18_next_int_m[4] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I3_G0N (.A(
        \state_RNI50LK1[0]_net_1 ), .B(average[3]), .Y(N326));
    AO13 un1_integ_0_0_ADD_26x26_fast_I48_Y (.A(LED_12[6]), .B(N353), 
        .C(\state_1[0]_net_1 ), .Y(N416));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I195_un1_Y (.A(N482), .B(N490), 
        .C(\state_1_RNIF5VI1[0]_net_1 ), .Y(I195_un1_Y));
    DFN1E0C0 \integ[3]  (.D(\un1_integ[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[3]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I252_Y (.A(I207_un1_Y), .B(
        ADD_26x26_fast_I207_Y_2), .C(ADD_26x26_fast_I252_Y_0), .Y(
        \un1_integ[22] ));
    DFN1E0C0 \integ[6]  (.D(\un1_integ[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[6]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_1 (.A(
        ADD_26x26_fast_I210_un1_Y_0), .B(N491), .C(
        ADD_26x26_fast_I210_Y_0), .Y(ADD_26x26_fast_I210_Y_1));
    NOR2B \state_RNIH8UP[0]  (.A(avg_new[4]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[4] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y (.A(N533), .B(I194_un1_Y), 
        .C(ADD_26x26_fast_I239_Y_0), .Y(\un1_integ[9] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I206_Y_0 (.A(N402), .B(N398), .Y(
        ADD_26x26_fast_I206_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I58_Y (.A(N338), .B(N342), .C(
        N341), .Y(N426));
    OA1 un1_integ_0_0_ADD_26x26_fast_I67_Y (.A(average[3]), .B(
        \state_RNI50LK1[0]_net_1 ), .C(N330), .Y(N435));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I253_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I253_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I64_Y (.A(N329), .B(N333), .C(
        N332), .Y(N432));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I204_un1_Y_0 (.A(N502), .B(N518)
        , .Y(ADD_26x26_fast_I204_un1_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I127_Y (.A(N401), .B(
        ADD_26x26_fast_I127_Y_0), .C(N458), .Y(N504));
    AO1 un1_integ_0_0_ADD_26x26_fast_I110_Y (.A(N432), .B(N429), .C(
        N428), .Y(N481));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I211_un1_Y_0 (.A(N462), .B(N470)
        , .C(N493), .Y(ADD_26x26_fast_I211_un1_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I90_Y (.A(N408), .B(N412), .Y(
        N461));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I233_Y (.A(
        \state_RNI50LK1[0]_net_1 ), .B(average[3]), .C(N491), .Y(
        \un1_integ[3] ));
    OA1A un1_integ_0_0_ADD_26x26_fast_I47_Y (.A(\state_1[0]_net_1 ), 
        .B(LED_12[7]), .C(N357), .Y(N415));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I119_Y (.A(N441), .B(N437), .Y(
        N490));
    AO1 un1_integ_0_0_ADD_26x26_fast_I70_Y (.A(N320), .B(N324), .C(
        N323), .Y(N438));
    NOR2B \state_1_RNIF0VM[0]  (.A(avg_new[11]), .B(\state_1[0]_net_1 )
        , .Y(\inf_abs0_m[11] ));
    DFN1E0C0 \integ[5]  (.D(\un1_integ[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[5]));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I182_un1_Y (.A(N462), .B(N470), 
        .C(N531), .Y(I182_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I161_Y (.A(N493), .B(N486), .C(
        N485), .Y(N539));
    OA1B un1_integ_0_0_ADD_26x26_fast_I44_Y (.A(LED_12[7]), .B(
        \integ[15]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N412));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I245_Y (.A(\state_1[0]_net_1 ), 
        .B(\integ[15]_net_1 ), .C(N637), .Y(\un1_integ[15] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I95_Y (.A(N417), .B(N413), .Y(
        N466));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y_0 (.A(
        \un18_next_int_m[9] ), .B(\inf_abs0_m[9] ), .C(LED_12[2]), .Y(
        ADD_26x26_fast_I239_Y_0));
    DFN1E0C0 \integ[2]  (.D(\un1_integ[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(average[2]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I135_Y (.A(N458), .B(N466), .Y(
        N512));
    OR2 un1_integ_0_0_ADD_26x26_fast_I88_Y (.A(N406), .B(N410), .Y(
        N459));
    AX1D un1_integ_0_0_ADD_26x26_fast_I247_Y (.A(I184_un1_Y), .B(
        ADD_26x26_fast_I212_Y_0), .C(ADD_26x26_fast_I247_Y_0), .Y(
        \un1_integ[17] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I143_Y (.A(N466), .B(N474), .Y(
        N520));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I57_Y (.A(N342), .B(N345), .Y(
        N425));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I186_un1_Y (.A(N535), .B(N520), 
        .Y(I186_un1_Y));
    DFN1E0C0 \integ[23]  (.D(\un1_integ[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[23]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I8_P0N (.A(\un1_next_int[8] ), .B(
        LED_12[1]), .Y(N342));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_2 (.A(N506), .B(N521), .C(
        ADD_26x26_fast_I206_Y_1), .Y(ADD_26x26_fast_I206_Y_2));
    AO1 un1_integ_0_0_ADD_26x26_fast_I54_Y (.A(N344), .B(N348), .C(
        N347), .Y(N422));
    NOR2A \state_RNIPSMQ[1]  (.A(\state[1]_net_1 ), .B(avg_old[7]), .Y(
        \un18_next_int_m[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I131_Y (.A(N454), .B(N462), .Y(
        N508));
    AX1D un1_integ_0_0_ADD_26x26_fast_I254_Y (.A(I205_un1_Y), .B(
        ADD_26x26_fast_I205_Y_3), .C(ADD_26x26_fast_I254_Y_0), .Y(
        \un1_integ[24] ));
    NOR2 \state_RNI9SUR[0]  (.A(\state[1]_net_1 ), .B(\state[0]_net_1 )
        , .Y(avg_done));
    NOR2A \state_RNI39TH[1]  (.A(\state[1]_net_1 ), .B(avg_old[10]), 
        .Y(\un18_next_int_m[10] ));
    DFN1E0C0 \integ[19]  (.D(\un1_integ[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[19]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I117_Y (.A(N439), .B(N435), .Y(
        N488));
    DFN1E0C0 \integ[17]  (.D(\un1_integ[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[17]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I33_Y (.A(\integ[21]_net_1 ), .B(
        \integ[20]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N401));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I255_Y_0 (.A(\integ[25]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I255_Y_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I127_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\integ[22]_net_1 ), .C(\state_1[0]_net_1 ), .Y(
        ADD_26x26_fast_I127_Y_0));
    DFN1E0C0 \integ[14]  (.D(\un1_integ[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_12[7]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I87_Y (.A(N405), .B(N409), .Y(
        N458));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y_0 (.A(average[2]), .B(
        \state_RNI3UKK1[0]_net_1 ), .Y(ADD_26x26_fast_I232_Y_0));
    NOR2A \state_RNILOMQ[1]  (.A(\state[1]_net_1 ), .B(avg_old[3]), .Y(
        \un18_next_int_m[3] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I84_Y (.A(N402), .B(N406), .Y(
        N455));
    AO1 un1_integ_0_0_ADD_26x26_fast_I154_Y (.A(N485), .B(N478), .C(
        N477), .Y(N531));
    OA1 un1_integ_0_0_ADD_26x26_fast_I11_G0N (.A(\un18_next_int_m[11] )
        , .B(\inf_abs0_m[11] ), .C(LED_12[4]), .Y(N350));
    AO1 un1_integ_0_0_ADD_26x26_fast_I140_Y (.A(N471), .B(N464), .C(
        N463), .Y(N517));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I149_Y (.A(N480), .B(N472), .Y(
        N526));
    AO1 un1_integ_0_0_ADD_26x26_fast_I158_Y (.A(N489), .B(N482), .C(
        N481), .Y(N535));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I249_Y_0 (.A(\integ[19]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I249_Y_0));
    DFN1E0C0 \integ[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done), .Q(\integ[25]_net_1 ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I247_Y_0 (.A(\integ[17]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I247_Y_0));
    NOR2A \un1_integ_0_0_LED_5[7]  (.A(LED_33[7]), .B(choose[2]), .Y(
        N_65));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y_0 (.A(\integ[0]_net_1 ), 
        .B(\state[1]_net_1 ), .Y(ADD_26x26_fast_I230_Y_0));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I242_Y (.A(\state[1]_net_1 ), .B(
        LED_12[5]), .C(N646), .Y(\un1_integ[12] ));
    DFN1E0C0 \integ[11]  (.D(\un1_integ[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(LED_12[4]));
    DFN1E0C0 \integ[16]  (.D(\un1_integ[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[16]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_1 (.A(
        ADD_26x26_fast_I211_un1_Y_0), .B(N532), .C(
        ADD_26x26_fast_I211_Y_0), .Y(ADD_26x26_fast_I211_Y_1));
    OR2 \state_RNI72LK1[0]  (.A(\inf_abs0_m[4] ), .B(
        \un18_next_int_m[4] ), .Y(\state_RNI72LK1[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I189_Y (.A(N524), .B(N539), .C(
        N523), .Y(N640));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I254_Y_0 (.A(\integ[24]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I254_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I163_Y (.A(I163_un1_Y), .B(N489), 
        .Y(N543));
    NOR2A \state_RNIQTMQ[1]  (.A(\state[1]_net_1 ), .B(avg_old[8]), .Y(
        \un18_next_int_m[8] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I96_Y (.A(N418), .B(N415), .C(
        N414), .Y(N467));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I207_un1_Y (.A(N524), .B(N508), 
        .C(N539), .Y(I207_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I2_G0N (.A(
        \state_RNI3UKK1[0]_net_1 ), .B(average[2]), .Y(N323));
    AO1 un1_integ_0_0_ADD_26x26_fast_I114_Y (.A(N436), .B(N433), .C(
        N432), .Y(N485));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I147_Y (.A(N470), .B(N478), .Y(
        N524));
    DFN1E0C0 \integ[9]  (.D(\un1_integ[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(LED_12[2]));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I235_Y (.A(
        ADD_26x26_fast_I235_Y_0), .B(N541), .Y(\un1_integ[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I212_Y_0 (.A(
        ADD_26x26_fast_I212_un1_Y_0), .B(N518), .C(N517), .Y(
        ADD_26x26_fast_I212_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I63_Y (.A(N333), .B(N336), .Y(
        N431));
    AO1 un1_integ_0_0_ADD_26x26_fast_I118_Y (.A(N440), .B(N437), .C(
        N436), .Y(N489));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I237_Y (.A(
        \state_RNID8LK1[0]_net_1 ), .B(LED_12[0]), .C(N537), .Y(
        \un1_integ[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I133_Y (.A(N456), .B(N464), .Y(
        N510));
    OA1B un1_integ_0_0_ADD_26x26_fast_I30_Y (.A(\integ[22]_net_1 ), .B(
        \integ[21]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N398));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I160_un1_Y (.A(N484), .B(N491), 
        .Y(I160_un1_Y));
    DFN1E0C0 \integ[22]  (.D(\un1_integ[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[22]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I43_Y (.A(\integ[15]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N411));
    DFN1E0C0 \integ[1]  (.D(\un1_integ[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(\integ[1]_net_1 ));
    MX2 \un1_integ_0_0_LED_1[7]  (.A(LED_12[7]), .B(LED_15[7]), .S(
        choose_0_0), .Y(N_104));
    AO1B un1_integ_0_0_ADD_26x26_fast_I35_Y (.A(\integ[20]_net_1 ), .B(
        \integ[19]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N403));
    OR2 \state_1_RNIF5VI1[0]  (.A(\inf_abs0_m[0] ), .B(
        \un18_next_int_m[0] ), .Y(\state_1_RNIF5VI1[0]_net_1 ));
    DFN1C0 \state_0[0]  (.D(\state_1_RNI4F701[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_0[0]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I53_Y (.A(N351), .B(N348), .Y(
        N421));
    OR2 un1_integ_0_0_ADD_26x26_fast_I160_Y (.A(I160_un1_Y), .B(N483), 
        .Y(N537));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I91_Y (.A(N413), .B(N409), .Y(
        N462));
    AX1D un1_integ_0_0_ADD_26x26_fast_I250_Y (.A(I178_un1_Y), .B(
        ADD_26x26_fast_I209_Y_1), .C(ADD_26x26_fast_I250_Y_0), .Y(
        \un1_integ[20] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I240_Y_0 (.A(LED_12[3]), .B(
        \state_1_RNIH8S81[0]_net_1 ), .Y(ADD_26x26_fast_I240_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_0 (.A(N467), .B(N460), .C(
        N459), .Y(ADD_26x26_fast_I210_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I71_Y (.A(N321), .B(N324), .Y(
        N439));
    DFN1E0C0 \integ[20]  (.D(\un1_integ[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[20]_net_1 ));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I244_Y (.A(\state_1[0]_net_1 ), 
        .B(LED_12[7]), .C(N640), .Y(\un1_integ[14] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_1 (.A(N461), .B(N454), .C(
        ADD_26x26_fast_I207_Y_0), .Y(ADD_26x26_fast_I207_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I106_Y (.A(N428), .B(N425), .C(
        N424), .Y(N477));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_1 (.A(
        ADD_26x26_fast_I208_un1_Y_0), .B(N541), .C(
        ADD_26x26_fast_I208_Y_0), .Y(ADD_26x26_fast_I208_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I102_Y (.A(N424), .B(N421), .C(
        N420), .Y(N473));
    NOR2B \state_RNIKBUP[0]  (.A(avg_new[7]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[7] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I251_Y (.A(I176_un1_Y), .B(
        ADD_26x26_fast_I208_Y_1), .C(ADD_26x26_fast_I251_Y_0), .Y(
        \un1_integ[21] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I121_un1_Y (.A(N441), .B(
        \state_1_RNIF5VI1[0]_net_1 ), .Y(I121_un1_Y));
    DFN1E0C0 \integ[18]  (.D(\un1_integ[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_done_0), .Q(\integ[18]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I4_P0N (.A(
        \state_RNI72LK1[0]_net_1 ), .B(average[4]), .Y(N330));
    NOR2A \un1_integ_0_0_LED_2[7]  (.A(LED_5[7]), .B(choose_0_0), .Y(
        N_41));
    AO1 un1_integ_0_0_ADD_26x26_fast_I144_Y (.A(N475), .B(N468), .C(
        N467), .Y(N521));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I83_Y (.A(N405), .B(N401), .Y(
        N454));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_0 (.A(N465), .B(N458), .C(
        N457), .Y(ADD_26x26_fast_I209_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I207_Y_0 (.A(N400), .B(N404), .Y(
        ADD_26x26_fast_I207_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I148_Y (.A(I148_un1_Y), .B(N471), 
        .Y(N525));
    MX2 \un1_integ_0_0_LED_3[7]  (.A(N_104), .B(N_41), .S(choose[1]), 
        .Y(N_49));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I60_Y (.A(N335), .B(
        \state_RNID8LK1[0]_net_1 ), .C(LED_12[0]), .Y(N428));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y (.A(
        ADD_26x26_fast_I232_Y_0), .B(N493), .Y(\un1_integ[2] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I204_Y_2 (.A(N398), .B(
        ADD_26x26_fast_I204_Y_0), .C(N455), .Y(ADD_26x26_fast_I204_Y_2)
        );
    DFN1C0 \state[1]  (.D(\state_RNO[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[1]_net_1 ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I9_G0N (.A(\un18_next_int_m[9] ), 
        .B(\inf_abs0_m[9] ), .C(LED_12[2]), .Y(N344));
    MX2 \un1_integ_0_0_LED_6[7]  (.A(N_57), .B(N_65), .S(choose[1]), 
        .Y(N_73));
    OA1B un1_integ_0_0_ADD_26x26_fast_I40_Y (.A(\integ[17]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N408));
    NOR2A \un1_integ_0_0_LED_4[6]  (.A(LED_FB[6]), .B(choose[2]), .Y(
        N_56));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I65_Y (.A(N333), .B(N330), .Y(
        N433));
    AO1 un1_integ_0_0_ADD_26x26_fast_I188_Y (.A(N522), .B(N537), .C(
        N521), .Y(N637));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I178_un1_Y (.A(N512), .B(N527), 
        .Y(I178_un1_Y));
    AO1B un1_integ_0_0_ADD_26x26_fast_I45_Y (.A(\integ[15]_net_1 ), .B(
        LED_12[7]), .C(\state_0[0]_net_1 ), .Y(N413));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I137_Y (.A(N460), .B(N468), .Y(
        N514));
    OR2 \state_RNIB6LK1[0]  (.A(\inf_abs0_m[6] ), .B(
        \un18_next_int_m[6] ), .Y(\state_RNIB6LK1[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I50_Y (.A(N350), .B(N354), .C(
        N353), .Y(N418));
    AO1 un1_integ_0_0_ADD_26x26_fast_I204_Y_3 (.A(N502), .B(N517), .C(
        ADD_26x26_fast_I204_Y_2), .Y(ADD_26x26_fast_I204_Y_3));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I74_un1_Y (.A(N318), .B(
        \state_1_RNIF5VI1[0]_net_1 ), .Y(I74_un1_Y));
    OA1B un1_integ_0_0_ADD_26x26_fast_I36_Y (.A(\integ[18]_net_1 ), .B(
        \integ[19]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N404));
    OR2 un1_integ_0_0_ADD_26x26_fast_I0_P0N (.A(\integ[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(N318));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I55_Y (.A(N345), .B(N348), .Y(
        N423));
    NOR2A \state_RNI4ATH[1]  (.A(\state[1]_net_1 ), .B(avg_old[11]), 
        .Y(\un18_next_int_m[11] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I205_un1_Y (.A(N535), .B(
        I195_un1_Y), .C(ADD_26x26_fast_I205_un1_Y_0), .Y(I205_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I163_un1_Y (.A(N490), .B(
        \state_1_RNIF5VI1[0]_net_1 ), .Y(I163_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_1 (.A(N452), .B(N459), .C(
        ADD_26x26_fast_I206_Y_0), .Y(ADD_26x26_fast_I206_Y_1));
    OA1 un1_integ_0_0_ADD_26x26_fast_I5_G0N (.A(\inf_abs0_m[5] ), .B(
        \un18_next_int_m[5] ), .C(average[5]), .Y(N332));
    OR2 \state_RNI50LK1[0]  (.A(\inf_abs0_m[3] ), .B(
        \un18_next_int_m[3] ), .Y(\state_RNI50LK1[0]_net_1 ));
    DFN1E0C0 \integ[7]  (.D(\un1_integ[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(LED_12[0]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_2 (.A(N508), .B(N523), .C(
        ADD_26x26_fast_I207_Y_1), .Y(ADD_26x26_fast_I207_Y_2));
    MX2 \un1_integ_0_0_LED_6[6]  (.A(N_56), .B(N_64), .S(choose[1]), 
        .Y(N_72));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I4_G0N (.A(
        \state_RNI72LK1[0]_net_1 ), .B(average[4]), .Y(N329));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I206_un1_Y_0 (.A(N506), .B(N522)
        , .Y(ADD_26x26_fast_I206_un1_Y_0));
    OR2 \state_RNIFALK1[0]  (.A(\un18_next_int_m[8] ), .B(
        \inf_abs0_m[8] ), .Y(\un1_next_int[8] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y (.A(
        ADD_26x26_fast_I234_Y_0), .B(N543), .Y(\un1_integ[4] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I205_Y_2 (.A(N400), .B(
        ADD_26x26_fast_I205_Y_0), .C(N457), .Y(ADD_26x26_fast_I205_Y_2)
        );
    NOR2B un1_integ_0_0_ADD_26x26_fast_I162_un1_Y (.A(N488), .B(N442), 
        .Y(I162_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I240_Y (.A(N531), .B(I193_un1_Y), 
        .C(ADD_26x26_fast_I240_Y_0), .Y(\un1_integ[10] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I156_Y (.A(N487), .B(N480), .C(
        N479), .Y(N533));
    DFN1E0C0 \integ[8]  (.D(\un1_integ[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(avg_done), .Q(LED_12[1]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I85_Y (.A(N407), .B(N403), .Y(
        N456));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I251_Y_0 (.A(\integ[21]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I251_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I152_Y (.A(I152_un1_Y), .B(N475), 
        .Y(N529));
    OR2 \state_RNID8LK1[0]  (.A(\inf_abs0_m[7] ), .B(
        \un18_next_int_m[7] ), .Y(\state_RNID8LK1[0]_net_1 ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I9_P0N (.A(\un18_next_int_m[9] ), 
        .B(\inf_abs0_m[9] ), .C(LED_12[2]), .Y(N345));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I208_un1_Y_0 (.A(N510), .B(N526)
        , .Y(ADD_26x26_fast_I208_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I191_Y (.A(N528), .B(N543), .C(
        N527), .Y(N646));
    AO1B un1_integ_0_0_ADD_26x26_fast_I31_Y (.A(\integ[21]_net_1 ), .B(
        \integ[22]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N399));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I206_un1_Y (.A(
        ADD_26x26_fast_I206_un1_Y_0), .B(N537), .Y(I206_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I235_Y_0 (.A(\inf_abs0_m[5] ), 
        .B(\un18_next_int_m[5] ), .C(average[5]), .Y(
        ADD_26x26_fast_I235_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I241_Y (.A(N529), .B(I192_un1_Y), 
        .C(ADD_26x26_fast_I241_Y_0), .Y(\un1_integ[11] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I11_P0N (.A(\un18_next_int_m[11] )
        , .B(\inf_abs0_m[11] ), .C(LED_12[4]), .Y(N351));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I105_Y (.A(N427), .B(N423), .Y(
        N476));
    AO1 un1_integ_0_0_ADD_26x26_fast_I213_Y_0 (.A(
        ADD_26x26_fast_I213_un1_Y_0), .B(N520), .C(N519), .Y(
        ADD_26x26_fast_I213_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I238_Y_0 (.A(LED_12[1]), .B(
        \un1_next_int[8] ), .Y(ADD_26x26_fast_I238_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I101_Y (.A(N419), .B(N423), .Y(
        N472));
    AO1 un1_integ_0_0_ADD_26x26_fast_I66_Y (.A(N326), .B(N330), .C(
        N329), .Y(N434));
    AX1D un1_integ_0_0_ADD_26x26_fast_I248_Y (.A(I182_un1_Y), .B(
        ADD_26x26_fast_I211_Y_1), .C(ADD_26x26_fast_I248_Y_0), .Y(
        \un1_integ[18] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I99_Y (.A(N417), .B(N421), .Y(
        N470));
    AO1 un1_integ_0_0_ADD_26x26_fast_I92_Y (.A(N414), .B(N411), .C(
        N410), .Y(N463));
    OR2 \state_RNI3UKK1[0]  (.A(\inf_abs0_m[2] ), .B(
        \un18_next_int_m[2] ), .Y(\state_RNI3UKK1[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I72_Y (.A(N317), .B(N321), .C(
        N320), .Y(N440));
    OR2A un1_integ_0_0_ADD_26x26_fast_I13_P0N (.A(\state_1[0]_net_1 ), 
        .B(LED_12[6]), .Y(N357));
    OA1B un1_integ_0_0_ADD_26x26_fast_I46_Y (.A(LED_12[7]), .B(
        LED_12[6]), .C(\state_0[0]_net_1 ), .Y(N414));
    NOR2B \state_1_RNITF8O[0]  (.A(avg_new[0]), .B(\state_1[0]_net_1 ), 
        .Y(\inf_abs0_m[0] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I116_Y (.A(N438), .B(N435), .C(
        N434), .Y(N487));
    AO1 un1_integ_0_0_ADD_26x26_fast_I112_Y (.A(N431), .B(N434), .C(
        N430), .Y(N483));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I8_G0N (.A(\un1_next_int[8] ), 
        .B(LED_12[1]), .Y(N341));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I213_un1_Y_0 (.A(N482), .B(N490)
        , .C(\state_1_RNIF5VI1[0]_net_1 ), .Y(
        ADD_26x26_fast_I213_un1_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y_0 (.A(average[4]), .B(
        \state_RNI72LK1[0]_net_1 ), .Y(ADD_26x26_fast_I234_Y_0));
    
endmodule


module error_sr_13s_5s(
       cur_vd,
       avg_new,
       avg_old,
       avg_enable_1,
       avg_enable_0,
       avg_enable,
       n_rst_c,
       clk_c
    );
input  [11:0] cur_vd;
output [11:0] avg_new;
output [11:0] avg_old;
input  avg_enable_1;
input  avg_enable_0;
input  avg_enable;
input  n_rst_c;
input  clk_c;

    wire \sr_3_[0]_net_1 , \sr_3_[1]_net_1 , \sr_3_[2]_net_1 , 
        \sr_3_[3]_net_1 , \sr_3_[4]_net_1 , \sr_3_[5]_net_1 , 
        \sr_3_[6]_net_1 , \sr_3_[7]_net_1 , \sr_3_[8]_net_1 , 
        \sr_3_[9]_net_1 , \sr_3_[10]_net_1 , \sr_3_[11]_net_1 , 
        \sr_2_[0]_net_1 , \sr_2_[1]_net_1 , \sr_2_[2]_net_1 , 
        \sr_2_[3]_net_1 , \sr_2_[4]_net_1 , \sr_2_[5]_net_1 , 
        \sr_2_[6]_net_1 , \sr_2_[7]_net_1 , \sr_2_[8]_net_1 , 
        \sr_2_[9]_net_1 , \sr_2_[10]_net_1 , \sr_2_[11]_net_1 , 
        \sr_1_[0]_net_1 , \sr_1_[1]_net_1 , \sr_1_[2]_net_1 , 
        \sr_1_[3]_net_1 , \sr_1_[4]_net_1 , \sr_1_[5]_net_1 , 
        \sr_1_[6]_net_1 , \sr_1_[7]_net_1 , \sr_1_[8]_net_1 , 
        \sr_1_[9]_net_1 , \sr_1_[10]_net_1 , \sr_1_[11]_net_1 , GND, 
        VCC;
    
    DFN1E1C0 \sr_1_[11]  (.D(avg_new[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(\sr_1_[11]_net_1 ));
    DFN1E1C0 \sr_3_[3]  (.D(\sr_2_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[3]_net_1 ));
    DFN1E1C0 \sr_4_[4]  (.D(\sr_3_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[4]));
    DFN1E1C0 \sr_0_[10]  (.D(cur_vd[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(avg_new[10]));
    DFN1E1C0 \sr_4_[8]  (.D(\sr_3_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[8]));
    DFN1E1C0 \sr_4_[0]  (.D(\sr_3_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[0]));
    DFN1E1C0 \sr_1_[2]  (.D(avg_new[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[2]_net_1 ));
    DFN1E1C0 \sr_0_[2]  (.D(cur_vd[2]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[2]));
    DFN1E1C0 \sr_2_[2]  (.D(\sr_1_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[2]_net_1 ));
    DFN1E1C0 \sr_0_[11]  (.D(cur_vd[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(avg_new[11]));
    DFN1E1C0 \sr_1_[3]  (.D(avg_new[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[3]_net_1 ));
    DFN1E1C0 \sr_0_[3]  (.D(cur_vd[3]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[3]));
    DFN1E1C0 \sr_1_[10]  (.D(avg_new[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_1), .Q(\sr_1_[10]_net_1 ));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \sr_4_[10]  (.D(\sr_3_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[10]));
    DFN1E1C0 \sr_3_[11]  (.D(\sr_2_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[11]_net_1 ));
    DFN1E1C0 \sr_2_[3]  (.D(\sr_1_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[3]_net_1 ));
    DFN1E1C0 \sr_3_[6]  (.D(\sr_2_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[6]_net_1 ));
    DFN1E1C0 \sr_3_[1]  (.D(\sr_2_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[1]_net_1 ));
    DFN1E1C0 \sr_4_[2]  (.D(\sr_3_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[2]));
    DFN1E1C0 \sr_1_[6]  (.D(avg_new[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[6]_net_1 ));
    DFN1E1C0 \sr_4_[3]  (.D(\sr_3_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[3]));
    DFN1E1C0 \sr_0_[6]  (.D(cur_vd[6]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[6]));
    DFN1E1C0 \sr_3_[9]  (.D(\sr_2_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[9]_net_1 ));
    DFN1E1C0 \sr_1_[1]  (.D(avg_new[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[1]_net_1 ));
    DFN1E1C0 \sr_0_[1]  (.D(cur_vd[1]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[1]));
    DFN1E1C0 \sr_2_[6]  (.D(\sr_1_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[6]_net_1 ));
    DFN1E1C0 \sr_2_[1]  (.D(\sr_1_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[1]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1C0 \sr_3_[5]  (.D(\sr_2_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[5]_net_1 ));
    DFN1E1C0 \sr_3_[7]  (.D(\sr_2_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[7]_net_1 ));
    DFN1E1C0 \sr_1_[9]  (.D(avg_new[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[9]_net_1 ));
    DFN1E1C0 \sr_0_[9]  (.D(cur_vd[9]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[9]));
    DFN1E1C0 \sr_2_[11]  (.D(\sr_1_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(\sr_2_[11]_net_1 ));
    DFN1E1C0 \sr_4_[6]  (.D(\sr_3_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[6]));
    DFN1E1C0 \sr_2_[9]  (.D(\sr_1_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[9]_net_1 ));
    DFN1E1C0 \sr_4_[11]  (.D(\sr_3_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(avg_old[11]));
    DFN1E1C0 \sr_4_[1]  (.D(\sr_3_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[1]));
    DFN1E1C0 \sr_3_[4]  (.D(\sr_2_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[4]_net_1 ));
    DFN1E1C0 \sr_1_[5]  (.D(avg_new[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[5]_net_1 ));
    DFN1E1C0 \sr_0_[5]  (.D(cur_vd[5]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[5]));
    DFN1E1C0 \sr_1_[7]  (.D(avg_new[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[7]_net_1 ));
    DFN1E1C0 \sr_0_[7]  (.D(cur_vd[7]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[7]));
    DFN1E1C0 \sr_3_[8]  (.D(\sr_2_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[8]_net_1 ));
    DFN1E1C0 \sr_3_[0]  (.D(\sr_2_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[0]_net_1 ));
    DFN1E1C0 \sr_2_[5]  (.D(\sr_1_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[5]_net_1 ));
    DFN1E1C0 \sr_2_[7]  (.D(\sr_1_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[7]_net_1 ));
    DFN1E1C0 \sr_4_[9]  (.D(\sr_3_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[9]));
    DFN1E1C0 \sr_1_[4]  (.D(avg_new[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[4]_net_1 ));
    DFN1E1C0 \sr_0_[4]  (.D(cur_vd[4]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[4]));
    DFN1E1C0 \sr_1_[8]  (.D(avg_new[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[8]_net_1 ));
    DFN1E1C0 \sr_1_[0]  (.D(avg_new[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[0]_net_1 ));
    DFN1E1C0 \sr_2_[4]  (.D(\sr_1_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[4]_net_1 ));
    DFN1E1C0 \sr_0_[8]  (.D(cur_vd[8]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable), .Q(avg_new[8]));
    DFN1E1C0 \sr_0_[0]  (.D(cur_vd[0]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[0]));
    DFN1E1C0 \sr_4_[5]  (.D(\sr_3_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[5]));
    DFN1E1C0 \sr_2_[8]  (.D(\sr_1_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[8]_net_1 ));
    DFN1E1C0 \sr_2_[0]  (.D(\sr_1_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[0]_net_1 ));
    DFN1E1C0 \sr_4_[7]  (.D(\sr_3_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[7]));
    DFN1E1C0 \sr_3_[10]  (.D(\sr_2_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[10]_net_1 ));
    DFN1E1C0 \sr_3_[2]  (.D(\sr_2_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[2]_net_1 ));
    DFN1E1C0 \sr_2_[10]  (.D(\sr_1_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(\sr_2_[10]_net_1 ));
    
endmodule


module error_sr_13s_64s(
       sr_old,
       sr_new,
       cur_error,
       sr_prev,
       sr_new_0_0,
       sr_new_1_0,
       int_enable,
       n_rst_c,
       clk_c
    );
output [12:0] sr_old;
output [12:0] sr_new;
input  [12:0] cur_error;
output [12:0] sr_prev;
output sr_new_0_0;
output sr_new_1_0;
input  int_enable;
input  n_rst_c;
input  clk_c;

    wire \sr_9_[0]_net_1 , \sr_8_[0]_net_1 , \sr_9_[1]_net_1 , 
        \sr_8_[1]_net_1 , \sr_9_[2]_net_1 , \sr_8_[2]_net_1 , 
        \sr_9_[3]_net_1 , \sr_8_[3]_net_1 , \sr_9_[4]_net_1 , 
        \sr_8_[4]_net_1 , \sr_9_[5]_net_1 , \sr_8_[5]_net_1 , 
        \sr_9_[6]_net_1 , \sr_8_[6]_net_1 , \sr_9_[7]_net_1 , 
        \sr_8_[7]_net_1 , \sr_9_[8]_net_1 , \sr_8_[8]_net_1 , 
        \sr_9_[9]_net_1 , \sr_8_[9]_net_1 , \sr_9_[10]_net_1 , 
        \sr_8_[10]_net_1 , \sr_9_[11]_net_1 , \sr_8_[11]_net_1 , 
        \sr_9_[12]_net_1 , \sr_8_[12]_net_1 , \sr_7_[0]_net_1 , 
        \sr_7_[1]_net_1 , \sr_7_[2]_net_1 , \sr_7_[3]_net_1 , 
        \sr_7_[4]_net_1 , \sr_7_[5]_net_1 , \sr_7_[6]_net_1 , 
        \sr_7_[7]_net_1 , \sr_7_[8]_net_1 , \sr_7_[9]_net_1 , 
        \sr_7_[10]_net_1 , \sr_7_[11]_net_1 , \sr_7_[12]_net_1 , 
        \sr_6_[0]_net_1 , \sr_6_[1]_net_1 , \sr_6_[2]_net_1 , 
        \sr_6_[3]_net_1 , \sr_6_[4]_net_1 , \sr_6_[5]_net_1 , 
        \sr_6_[6]_net_1 , \sr_6_[7]_net_1 , \sr_6_[8]_net_1 , 
        \sr_6_[9]_net_1 , \sr_6_[10]_net_1 , \sr_6_[11]_net_1 , 
        \sr_6_[12]_net_1 , \sr_5_[0]_net_1 , \sr_5_[1]_net_1 , 
        \sr_5_[2]_net_1 , \sr_5_[3]_net_1 , \sr_5_[4]_net_1 , 
        \sr_5_[5]_net_1 , \sr_5_[6]_net_1 , \sr_5_[7]_net_1 , 
        \sr_5_[8]_net_1 , \sr_5_[9]_net_1 , \sr_5_[10]_net_1 , 
        \sr_5_[11]_net_1 , \sr_5_[12]_net_1 , \sr_4_[0]_net_1 , 
        \sr_4_[1]_net_1 , \sr_4_[2]_net_1 , \sr_4_[3]_net_1 , 
        \sr_4_[4]_net_1 , \sr_4_[5]_net_1 , \sr_4_[6]_net_1 , 
        \sr_4_[7]_net_1 , \sr_4_[8]_net_1 , \sr_4_[9]_net_1 , 
        \sr_4_[10]_net_1 , \sr_4_[11]_net_1 , \sr_4_[12]_net_1 , 
        \sr_3_[0]_net_1 , \sr_3_[1]_net_1 , \sr_3_[2]_net_1 , 
        \sr_3_[3]_net_1 , \sr_3_[4]_net_1 , \sr_3_[5]_net_1 , 
        \sr_3_[6]_net_1 , \sr_3_[7]_net_1 , \sr_3_[8]_net_1 , 
        \sr_3_[9]_net_1 , \sr_3_[10]_net_1 , \sr_3_[11]_net_1 , 
        \sr_3_[12]_net_1 , \sr_2_[0]_net_1 , \sr_2_[1]_net_1 , 
        \sr_2_[2]_net_1 , \sr_2_[3]_net_1 , \sr_2_[4]_net_1 , 
        \sr_2_[5]_net_1 , \sr_2_[6]_net_1 , \sr_2_[7]_net_1 , 
        \sr_2_[8]_net_1 , \sr_2_[9]_net_1 , \sr_2_[10]_net_1 , 
        \sr_2_[11]_net_1 , \sr_2_[12]_net_1 , \sr_24_[0]_net_1 , 
        \sr_23_[0]_net_1 , \sr_24_[1]_net_1 , \sr_23_[1]_net_1 , 
        \sr_24_[2]_net_1 , \sr_23_[2]_net_1 , \sr_24_[3]_net_1 , 
        \sr_23_[3]_net_1 , \sr_24_[4]_net_1 , \sr_23_[4]_net_1 , 
        \sr_24_[5]_net_1 , \sr_23_[5]_net_1 , \sr_24_[6]_net_1 , 
        \sr_23_[6]_net_1 , \sr_24_[7]_net_1 , \sr_23_[7]_net_1 , 
        \sr_24_[8]_net_1 , \sr_23_[8]_net_1 , \sr_24_[9]_net_1 , 
        \sr_23_[9]_net_1 , \sr_24_[10]_net_1 , \sr_23_[10]_net_1 , 
        \sr_24_[11]_net_1 , \sr_23_[11]_net_1 , \sr_24_[12]_net_1 , 
        \sr_23_[12]_net_1 , \sr_22_[0]_net_1 , \sr_22_[1]_net_1 , 
        \sr_22_[2]_net_1 , \sr_22_[3]_net_1 , \sr_22_[4]_net_1 , 
        \sr_22_[5]_net_1 , \sr_22_[6]_net_1 , \sr_22_[7]_net_1 , 
        \sr_22_[8]_net_1 , \sr_22_[9]_net_1 , \sr_22_[10]_net_1 , 
        \sr_22_[11]_net_1 , \sr_22_[12]_net_1 , \sr_21_[0]_net_1 , 
        \sr_21_[1]_net_1 , \sr_21_[2]_net_1 , \sr_21_[3]_net_1 , 
        \sr_21_[4]_net_1 , \sr_21_[5]_net_1 , \sr_21_[6]_net_1 , 
        \sr_21_[7]_net_1 , \sr_21_[8]_net_1 , \sr_21_[9]_net_1 , 
        \sr_21_[10]_net_1 , \sr_21_[11]_net_1 , \sr_21_[12]_net_1 , 
        \sr_20_[0]_net_1 , \sr_20_[1]_net_1 , \sr_20_[2]_net_1 , 
        \sr_20_[3]_net_1 , \sr_20_[4]_net_1 , \sr_20_[5]_net_1 , 
        \sr_20_[6]_net_1 , \sr_20_[7]_net_1 , \sr_20_[8]_net_1 , 
        \sr_20_[9]_net_1 , \sr_20_[10]_net_1 , \sr_20_[11]_net_1 , 
        \sr_20_[12]_net_1 , \sr_19_[0]_net_1 , \sr_19_[1]_net_1 , 
        \sr_19_[2]_net_1 , \sr_19_[3]_net_1 , \sr_19_[4]_net_1 , 
        \sr_19_[5]_net_1 , \sr_19_[6]_net_1 , \sr_19_[7]_net_1 , 
        \sr_19_[8]_net_1 , \sr_19_[9]_net_1 , \sr_19_[10]_net_1 , 
        \sr_19_[11]_net_1 , \sr_19_[12]_net_1 , \sr_18_[0]_net_1 , 
        \sr_18_[1]_net_1 , \sr_18_[2]_net_1 , \sr_18_[3]_net_1 , 
        \sr_18_[4]_net_1 , \sr_18_[5]_net_1 , \sr_18_[6]_net_1 , 
        \sr_18_[7]_net_1 , \sr_18_[8]_net_1 , \sr_18_[9]_net_1 , 
        \sr_18_[10]_net_1 , \sr_18_[11]_net_1 , \sr_18_[12]_net_1 , 
        \sr_17_[0]_net_1 , \sr_17_[1]_net_1 , \sr_17_[2]_net_1 , 
        \sr_17_[3]_net_1 , \sr_17_[4]_net_1 , \sr_17_[5]_net_1 , 
        \sr_17_[6]_net_1 , \sr_17_[7]_net_1 , \sr_17_[8]_net_1 , 
        \sr_17_[9]_net_1 , \sr_17_[10]_net_1 , \sr_17_[11]_net_1 , 
        \sr_17_[12]_net_1 , \sr_16_[0]_net_1 , \sr_16_[1]_net_1 , 
        \sr_16_[2]_net_1 , \sr_16_[3]_net_1 , \sr_16_[4]_net_1 , 
        \sr_16_[5]_net_1 , \sr_16_[6]_net_1 , \sr_16_[7]_net_1 , 
        \sr_16_[8]_net_1 , \sr_16_[9]_net_1 , \sr_16_[10]_net_1 , 
        \sr_16_[11]_net_1 , \sr_16_[12]_net_1 , \sr_15_[0]_net_1 , 
        \sr_15_[1]_net_1 , \sr_15_[2]_net_1 , \sr_15_[3]_net_1 , 
        \sr_15_[4]_net_1 , \sr_15_[5]_net_1 , \sr_15_[6]_net_1 , 
        \sr_15_[7]_net_1 , \sr_15_[8]_net_1 , \sr_15_[9]_net_1 , 
        \sr_15_[10]_net_1 , \sr_15_[11]_net_1 , \sr_15_[12]_net_1 , 
        \sr_14_[0]_net_1 , \sr_14_[1]_net_1 , \sr_14_[2]_net_1 , 
        \sr_14_[3]_net_1 , \sr_14_[4]_net_1 , \sr_14_[5]_net_1 , 
        \sr_14_[6]_net_1 , \sr_14_[7]_net_1 , \sr_14_[8]_net_1 , 
        \sr_14_[9]_net_1 , \sr_14_[10]_net_1 , \sr_14_[11]_net_1 , 
        \sr_14_[12]_net_1 , \sr_13_[0]_net_1 , \sr_13_[1]_net_1 , 
        \sr_13_[2]_net_1 , \sr_13_[3]_net_1 , \sr_13_[4]_net_1 , 
        \sr_13_[5]_net_1 , \sr_13_[6]_net_1 , \sr_13_[7]_net_1 , 
        \sr_13_[8]_net_1 , \sr_13_[9]_net_1 , \sr_13_[10]_net_1 , 
        \sr_13_[11]_net_1 , \sr_13_[12]_net_1 , \sr_12_[0]_net_1 , 
        \sr_12_[1]_net_1 , \sr_12_[2]_net_1 , \sr_12_[3]_net_1 , 
        \sr_12_[4]_net_1 , \sr_12_[5]_net_1 , \sr_12_[6]_net_1 , 
        \sr_12_[7]_net_1 , \sr_12_[8]_net_1 , \sr_12_[9]_net_1 , 
        \sr_12_[10]_net_1 , \sr_12_[11]_net_1 , \sr_12_[12]_net_1 , 
        \sr_11_[0]_net_1 , \sr_11_[1]_net_1 , \sr_11_[2]_net_1 , 
        \sr_11_[3]_net_1 , \sr_11_[4]_net_1 , \sr_11_[5]_net_1 , 
        \sr_11_[6]_net_1 , \sr_11_[7]_net_1 , \sr_11_[8]_net_1 , 
        \sr_11_[9]_net_1 , \sr_11_[10]_net_1 , \sr_11_[11]_net_1 , 
        \sr_11_[12]_net_1 , \sr_10_[0]_net_1 , \sr_10_[1]_net_1 , 
        \sr_10_[2]_net_1 , \sr_10_[3]_net_1 , \sr_10_[4]_net_1 , 
        \sr_10_[5]_net_1 , \sr_10_[6]_net_1 , \sr_10_[7]_net_1 , 
        \sr_10_[8]_net_1 , \sr_10_[9]_net_1 , \sr_10_[10]_net_1 , 
        \sr_10_[11]_net_1 , \sr_10_[12]_net_1 , \sr_39_[0]_net_1 , 
        \sr_38_[0]_net_1 , \sr_39_[1]_net_1 , \sr_38_[1]_net_1 , 
        \sr_39_[2]_net_1 , \sr_38_[2]_net_1 , \sr_39_[3]_net_1 , 
        \sr_38_[3]_net_1 , \sr_39_[4]_net_1 , \sr_38_[4]_net_1 , 
        \sr_39_[5]_net_1 , \sr_38_[5]_net_1 , \sr_39_[6]_net_1 , 
        \sr_38_[6]_net_1 , \sr_39_[7]_net_1 , \sr_38_[7]_net_1 , 
        \sr_39_[8]_net_1 , \sr_38_[8]_net_1 , \sr_39_[9]_net_1 , 
        \sr_38_[9]_net_1 , \sr_39_[10]_net_1 , \sr_38_[10]_net_1 , 
        \sr_39_[11]_net_1 , \sr_38_[11]_net_1 , \sr_39_[12]_net_1 , 
        \sr_38_[12]_net_1 , \sr_37_[0]_net_1 , \sr_37_[1]_net_1 , 
        \sr_37_[2]_net_1 , \sr_37_[3]_net_1 , \sr_37_[4]_net_1 , 
        \sr_37_[5]_net_1 , \sr_37_[6]_net_1 , \sr_37_[7]_net_1 , 
        \sr_37_[8]_net_1 , \sr_37_[9]_net_1 , \sr_37_[10]_net_1 , 
        \sr_37_[11]_net_1 , \sr_37_[12]_net_1 , \sr_36_[0]_net_1 , 
        \sr_36_[1]_net_1 , \sr_36_[2]_net_1 , \sr_36_[3]_net_1 , 
        \sr_36_[4]_net_1 , \sr_36_[5]_net_1 , \sr_36_[6]_net_1 , 
        \sr_36_[7]_net_1 , \sr_36_[8]_net_1 , \sr_36_[9]_net_1 , 
        \sr_36_[10]_net_1 , \sr_36_[11]_net_1 , \sr_36_[12]_net_1 , 
        \sr_35_[0]_net_1 , \sr_35_[1]_net_1 , \sr_35_[2]_net_1 , 
        \sr_35_[3]_net_1 , \sr_35_[4]_net_1 , \sr_35_[5]_net_1 , 
        \sr_35_[6]_net_1 , \sr_35_[7]_net_1 , \sr_35_[8]_net_1 , 
        \sr_35_[9]_net_1 , \sr_35_[10]_net_1 , \sr_35_[11]_net_1 , 
        \sr_35_[12]_net_1 , \sr_34_[0]_net_1 , \sr_34_[1]_net_1 , 
        \sr_34_[2]_net_1 , \sr_34_[3]_net_1 , \sr_34_[4]_net_1 , 
        \sr_34_[5]_net_1 , \sr_34_[6]_net_1 , \sr_34_[7]_net_1 , 
        \sr_34_[8]_net_1 , \sr_34_[9]_net_1 , \sr_34_[10]_net_1 , 
        \sr_34_[11]_net_1 , \sr_34_[12]_net_1 , \sr_33_[0]_net_1 , 
        \sr_33_[1]_net_1 , \sr_33_[2]_net_1 , \sr_33_[3]_net_1 , 
        \sr_33_[4]_net_1 , \sr_33_[5]_net_1 , \sr_33_[6]_net_1 , 
        \sr_33_[7]_net_1 , \sr_33_[8]_net_1 , \sr_33_[9]_net_1 , 
        \sr_33_[10]_net_1 , \sr_33_[11]_net_1 , \sr_33_[12]_net_1 , 
        \sr_32_[0]_net_1 , \sr_32_[1]_net_1 , \sr_32_[2]_net_1 , 
        \sr_32_[3]_net_1 , \sr_32_[4]_net_1 , \sr_32_[5]_net_1 , 
        \sr_32_[6]_net_1 , \sr_32_[7]_net_1 , \sr_32_[8]_net_1 , 
        \sr_32_[9]_net_1 , \sr_32_[10]_net_1 , \sr_32_[11]_net_1 , 
        \sr_32_[12]_net_1 , \sr_31_[0]_net_1 , \sr_31_[1]_net_1 , 
        \sr_31_[2]_net_1 , \sr_31_[3]_net_1 , \sr_31_[4]_net_1 , 
        \sr_31_[5]_net_1 , \sr_31_[6]_net_1 , \sr_31_[7]_net_1 , 
        \sr_31_[8]_net_1 , \sr_31_[9]_net_1 , \sr_31_[10]_net_1 , 
        \sr_31_[11]_net_1 , \sr_31_[12]_net_1 , \sr_30_[0]_net_1 , 
        \sr_30_[1]_net_1 , \sr_30_[2]_net_1 , \sr_30_[3]_net_1 , 
        \sr_30_[4]_net_1 , \sr_30_[5]_net_1 , \sr_30_[6]_net_1 , 
        \sr_30_[7]_net_1 , \sr_30_[8]_net_1 , \sr_30_[9]_net_1 , 
        \sr_30_[10]_net_1 , \sr_30_[11]_net_1 , \sr_30_[12]_net_1 , 
        \sr_29_[0]_net_1 , \sr_29_[1]_net_1 , \sr_29_[2]_net_1 , 
        \sr_29_[3]_net_1 , \sr_29_[4]_net_1 , \sr_29_[5]_net_1 , 
        \sr_29_[6]_net_1 , \sr_29_[7]_net_1 , \sr_29_[8]_net_1 , 
        \sr_29_[9]_net_1 , \sr_29_[10]_net_1 , \sr_29_[11]_net_1 , 
        \sr_29_[12]_net_1 , \sr_28_[0]_net_1 , \sr_28_[1]_net_1 , 
        \sr_28_[2]_net_1 , \sr_28_[3]_net_1 , \sr_28_[4]_net_1 , 
        \sr_28_[5]_net_1 , \sr_28_[6]_net_1 , \sr_28_[7]_net_1 , 
        \sr_28_[8]_net_1 , \sr_28_[9]_net_1 , \sr_28_[10]_net_1 , 
        \sr_28_[11]_net_1 , \sr_28_[12]_net_1 , \sr_27_[0]_net_1 , 
        \sr_27_[1]_net_1 , \sr_27_[2]_net_1 , \sr_27_[3]_net_1 , 
        \sr_27_[4]_net_1 , \sr_27_[5]_net_1 , \sr_27_[6]_net_1 , 
        \sr_27_[7]_net_1 , \sr_27_[8]_net_1 , \sr_27_[9]_net_1 , 
        \sr_27_[10]_net_1 , \sr_27_[11]_net_1 , \sr_27_[12]_net_1 , 
        \sr_26_[0]_net_1 , \sr_26_[1]_net_1 , \sr_26_[2]_net_1 , 
        \sr_26_[3]_net_1 , \sr_26_[4]_net_1 , \sr_26_[5]_net_1 , 
        \sr_26_[6]_net_1 , \sr_26_[7]_net_1 , \sr_26_[8]_net_1 , 
        \sr_26_[9]_net_1 , \sr_26_[10]_net_1 , \sr_26_[11]_net_1 , 
        \sr_26_[12]_net_1 , \sr_25_[0]_net_1 , \sr_25_[1]_net_1 , 
        \sr_25_[2]_net_1 , \sr_25_[3]_net_1 , \sr_25_[4]_net_1 , 
        \sr_25_[5]_net_1 , \sr_25_[6]_net_1 , \sr_25_[7]_net_1 , 
        \sr_25_[8]_net_1 , \sr_25_[9]_net_1 , \sr_25_[10]_net_1 , 
        \sr_25_[11]_net_1 , \sr_25_[12]_net_1 , \sr_54_[0]_net_1 , 
        \sr_53_[0]_net_1 , \sr_54_[1]_net_1 , \sr_53_[1]_net_1 , 
        \sr_54_[2]_net_1 , \sr_53_[2]_net_1 , \sr_54_[3]_net_1 , 
        \sr_53_[3]_net_1 , \sr_54_[4]_net_1 , \sr_53_[4]_net_1 , 
        \sr_54_[5]_net_1 , \sr_53_[5]_net_1 , \sr_54_[6]_net_1 , 
        \sr_53_[6]_net_1 , \sr_54_[7]_net_1 , \sr_53_[7]_net_1 , 
        \sr_54_[8]_net_1 , \sr_53_[8]_net_1 , \sr_54_[9]_net_1 , 
        \sr_53_[9]_net_1 , \sr_54_[10]_net_1 , \sr_53_[10]_net_1 , 
        \sr_54_[11]_net_1 , \sr_53_[11]_net_1 , \sr_54_[12]_net_1 , 
        \sr_53_[12]_net_1 , \sr_52_[0]_net_1 , \sr_52_[1]_net_1 , 
        \sr_52_[2]_net_1 , \sr_52_[3]_net_1 , \sr_52_[4]_net_1 , 
        \sr_52_[5]_net_1 , \sr_52_[6]_net_1 , \sr_52_[7]_net_1 , 
        \sr_52_[8]_net_1 , \sr_52_[9]_net_1 , \sr_52_[10]_net_1 , 
        \sr_52_[11]_net_1 , \sr_52_[12]_net_1 , \sr_51_[0]_net_1 , 
        \sr_51_[1]_net_1 , \sr_51_[2]_net_1 , \sr_51_[3]_net_1 , 
        \sr_51_[4]_net_1 , \sr_51_[5]_net_1 , \sr_51_[6]_net_1 , 
        \sr_51_[7]_net_1 , \sr_51_[8]_net_1 , \sr_51_[9]_net_1 , 
        \sr_51_[10]_net_1 , \sr_51_[11]_net_1 , \sr_51_[12]_net_1 , 
        \sr_50_[0]_net_1 , \sr_50_[1]_net_1 , \sr_50_[2]_net_1 , 
        \sr_50_[3]_net_1 , \sr_50_[4]_net_1 , \sr_50_[5]_net_1 , 
        \sr_50_[6]_net_1 , \sr_50_[7]_net_1 , \sr_50_[8]_net_1 , 
        \sr_50_[9]_net_1 , \sr_50_[10]_net_1 , \sr_50_[11]_net_1 , 
        \sr_50_[12]_net_1 , \sr_49_[0]_net_1 , \sr_49_[1]_net_1 , 
        \sr_49_[2]_net_1 , \sr_49_[3]_net_1 , \sr_49_[4]_net_1 , 
        \sr_49_[5]_net_1 , \sr_49_[6]_net_1 , \sr_49_[7]_net_1 , 
        \sr_49_[8]_net_1 , \sr_49_[9]_net_1 , \sr_49_[10]_net_1 , 
        \sr_49_[11]_net_1 , \sr_49_[12]_net_1 , \sr_48_[0]_net_1 , 
        \sr_48_[1]_net_1 , \sr_48_[2]_net_1 , \sr_48_[3]_net_1 , 
        \sr_48_[4]_net_1 , \sr_48_[5]_net_1 , \sr_48_[6]_net_1 , 
        \sr_48_[7]_net_1 , \sr_48_[8]_net_1 , \sr_48_[9]_net_1 , 
        \sr_48_[10]_net_1 , \sr_48_[11]_net_1 , \sr_48_[12]_net_1 , 
        \sr_47_[0]_net_1 , \sr_47_[1]_net_1 , \sr_47_[2]_net_1 , 
        \sr_47_[3]_net_1 , \sr_47_[4]_net_1 , \sr_47_[5]_net_1 , 
        \sr_47_[6]_net_1 , \sr_47_[7]_net_1 , \sr_47_[8]_net_1 , 
        \sr_47_[9]_net_1 , \sr_47_[10]_net_1 , \sr_47_[11]_net_1 , 
        \sr_47_[12]_net_1 , \sr_46_[0]_net_1 , \sr_46_[1]_net_1 , 
        \sr_46_[2]_net_1 , \sr_46_[3]_net_1 , \sr_46_[4]_net_1 , 
        \sr_46_[5]_net_1 , \sr_46_[6]_net_1 , \sr_46_[7]_net_1 , 
        \sr_46_[8]_net_1 , \sr_46_[9]_net_1 , \sr_46_[10]_net_1 , 
        \sr_46_[11]_net_1 , \sr_46_[12]_net_1 , \sr_45_[0]_net_1 , 
        \sr_45_[1]_net_1 , \sr_45_[2]_net_1 , \sr_45_[3]_net_1 , 
        \sr_45_[4]_net_1 , \sr_45_[5]_net_1 , \sr_45_[6]_net_1 , 
        \sr_45_[7]_net_1 , \sr_45_[8]_net_1 , \sr_45_[9]_net_1 , 
        \sr_45_[10]_net_1 , \sr_45_[11]_net_1 , \sr_45_[12]_net_1 , 
        \sr_44_[0]_net_1 , \sr_44_[1]_net_1 , \sr_44_[2]_net_1 , 
        \sr_44_[3]_net_1 , \sr_44_[4]_net_1 , \sr_44_[5]_net_1 , 
        \sr_44_[6]_net_1 , \sr_44_[7]_net_1 , \sr_44_[8]_net_1 , 
        \sr_44_[9]_net_1 , \sr_44_[10]_net_1 , \sr_44_[11]_net_1 , 
        \sr_44_[12]_net_1 , \sr_43_[0]_net_1 , \sr_43_[1]_net_1 , 
        \sr_43_[2]_net_1 , \sr_43_[3]_net_1 , \sr_43_[4]_net_1 , 
        \sr_43_[5]_net_1 , \sr_43_[6]_net_1 , \sr_43_[7]_net_1 , 
        \sr_43_[8]_net_1 , \sr_43_[9]_net_1 , \sr_43_[10]_net_1 , 
        \sr_43_[11]_net_1 , \sr_43_[12]_net_1 , \sr_42_[0]_net_1 , 
        \sr_42_[1]_net_1 , \sr_42_[2]_net_1 , \sr_42_[3]_net_1 , 
        \sr_42_[4]_net_1 , \sr_42_[5]_net_1 , \sr_42_[6]_net_1 , 
        \sr_42_[7]_net_1 , \sr_42_[8]_net_1 , \sr_42_[9]_net_1 , 
        \sr_42_[10]_net_1 , \sr_42_[11]_net_1 , \sr_42_[12]_net_1 , 
        \sr_41_[0]_net_1 , \sr_41_[1]_net_1 , \sr_41_[2]_net_1 , 
        \sr_41_[3]_net_1 , \sr_41_[4]_net_1 , \sr_41_[5]_net_1 , 
        \sr_41_[6]_net_1 , \sr_41_[7]_net_1 , \sr_41_[8]_net_1 , 
        \sr_41_[9]_net_1 , \sr_41_[10]_net_1 , \sr_41_[11]_net_1 , 
        \sr_41_[12]_net_1 , \sr_40_[0]_net_1 , \sr_40_[1]_net_1 , 
        \sr_40_[2]_net_1 , \sr_40_[3]_net_1 , \sr_40_[4]_net_1 , 
        \sr_40_[5]_net_1 , \sr_40_[6]_net_1 , \sr_40_[7]_net_1 , 
        \sr_40_[8]_net_1 , \sr_40_[9]_net_1 , \sr_40_[10]_net_1 , 
        \sr_40_[11]_net_1 , \sr_40_[12]_net_1 , \sr_62_[0]_net_1 , 
        \sr_62_[1]_net_1 , \sr_62_[2]_net_1 , \sr_62_[3]_net_1 , 
        \sr_62_[4]_net_1 , \sr_62_[5]_net_1 , \sr_62_[6]_net_1 , 
        \sr_62_[7]_net_1 , \sr_62_[8]_net_1 , \sr_62_[9]_net_1 , 
        \sr_62_[10]_net_1 , \sr_62_[11]_net_1 , \sr_62_[12]_net_1 , 
        \sr_61_[0]_net_1 , \sr_61_[1]_net_1 , \sr_61_[2]_net_1 , 
        \sr_61_[3]_net_1 , \sr_61_[4]_net_1 , \sr_61_[5]_net_1 , 
        \sr_61_[6]_net_1 , \sr_61_[7]_net_1 , \sr_61_[8]_net_1 , 
        \sr_61_[9]_net_1 , \sr_61_[10]_net_1 , \sr_61_[11]_net_1 , 
        \sr_61_[12]_net_1 , \sr_60_[0]_net_1 , \sr_60_[1]_net_1 , 
        \sr_60_[2]_net_1 , \sr_60_[3]_net_1 , \sr_60_[4]_net_1 , 
        \sr_60_[5]_net_1 , \sr_60_[6]_net_1 , \sr_60_[7]_net_1 , 
        \sr_60_[8]_net_1 , \sr_60_[9]_net_1 , \sr_60_[10]_net_1 , 
        \sr_60_[11]_net_1 , \sr_60_[12]_net_1 , \sr_59_[0]_net_1 , 
        \sr_59_[1]_net_1 , \sr_59_[2]_net_1 , \sr_59_[3]_net_1 , 
        \sr_59_[4]_net_1 , \sr_59_[5]_net_1 , \sr_59_[6]_net_1 , 
        \sr_59_[7]_net_1 , \sr_59_[8]_net_1 , \sr_59_[9]_net_1 , 
        \sr_59_[10]_net_1 , \sr_59_[11]_net_1 , \sr_59_[12]_net_1 , 
        \sr_58_[0]_net_1 , \sr_58_[1]_net_1 , \sr_58_[2]_net_1 , 
        \sr_58_[3]_net_1 , \sr_58_[4]_net_1 , \sr_58_[5]_net_1 , 
        \sr_58_[6]_net_1 , \sr_58_[7]_net_1 , \sr_58_[8]_net_1 , 
        \sr_58_[9]_net_1 , \sr_58_[10]_net_1 , \sr_58_[11]_net_1 , 
        \sr_58_[12]_net_1 , \sr_57_[0]_net_1 , \sr_57_[1]_net_1 , 
        \sr_57_[2]_net_1 , \sr_57_[3]_net_1 , \sr_57_[4]_net_1 , 
        \sr_57_[5]_net_1 , \sr_57_[6]_net_1 , \sr_57_[7]_net_1 , 
        \sr_57_[8]_net_1 , \sr_57_[9]_net_1 , \sr_57_[10]_net_1 , 
        \sr_57_[11]_net_1 , \sr_57_[12]_net_1 , \sr_56_[0]_net_1 , 
        \sr_56_[1]_net_1 , \sr_56_[2]_net_1 , \sr_56_[3]_net_1 , 
        \sr_56_[4]_net_1 , \sr_56_[5]_net_1 , \sr_56_[6]_net_1 , 
        \sr_56_[7]_net_1 , \sr_56_[8]_net_1 , \sr_56_[9]_net_1 , 
        \sr_56_[10]_net_1 , \sr_56_[11]_net_1 , \sr_56_[12]_net_1 , 
        \sr_55_[0]_net_1 , \sr_55_[1]_net_1 , \sr_55_[2]_net_1 , 
        \sr_55_[3]_net_1 , \sr_55_[4]_net_1 , \sr_55_[5]_net_1 , 
        \sr_55_[6]_net_1 , \sr_55_[7]_net_1 , \sr_55_[8]_net_1 , 
        \sr_55_[9]_net_1 , \sr_55_[10]_net_1 , \sr_55_[11]_net_1 , 
        \sr_55_[12]_net_1 , GND, VCC;
    
    DFN1E1C0 \sr_41_[5]  (.D(\sr_40_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[5]_net_1 ));
    DFN1E1C0 \sr_15_[3]  (.D(\sr_14_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[3]_net_1 ));
    DFN1E1C0 \sr_36_[5]  (.D(\sr_35_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[5]_net_1 ));
    DFN1E1C0 \sr_57_[5]  (.D(\sr_56_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[5]_net_1 ));
    DFN1E1C0 \sr_45_[11]  (.D(\sr_44_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[11]_net_1 ));
    DFN1E1C0 \sr_39_[6]  (.D(\sr_38_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[6]_net_1 ));
    DFN1E1C0 \sr_36_[4]  (.D(\sr_35_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[4]_net_1 ));
    DFN1E1C0 \sr_42_[4]  (.D(\sr_41_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[4]_net_1 ));
    DFN1E1C0 \sr_9_[3]  (.D(\sr_8_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[3]_net_1 ));
    DFN1E1C0 \sr_6_[4]  (.D(\sr_5_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[4]_net_1 ));
    DFN1E1C0 \sr_32_[3]  (.D(\sr_31_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[3]_net_1 ));
    DFN1E1C0 \sr_52_[6]  (.D(\sr_51_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[6]_net_1 ));
    DFN1E1C0 \sr_21_[9]  (.D(\sr_20_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[9]_net_1 ));
    DFN1E1C0 \sr_47_[12]  (.D(\sr_46_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[12]_net_1 ));
    DFN1E1C0 \sr_22_[4]  (.D(\sr_21_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[4]_net_1 ));
    DFN1E1C0 \sr_10_[1]  (.D(\sr_9_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[1]_net_1 ));
    DFN1E1C0 \sr_5_[4]  (.D(\sr_4_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[4]_net_1 ));
    DFN1E1C0 \sr_62_[6]  (.D(\sr_61_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[6]_net_1 ));
    DFN1E1C0 \sr_58_[2]  (.D(\sr_57_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[2]_net_1 ));
    DFN1E1C0 \sr_55_[0]  (.D(\sr_54_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[0]_net_1 ));
    DFN1E1C0 \sr_27_[3]  (.D(\sr_26_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[3]_net_1 ));
    DFN1E1C0 \sr_21_[1]  (.D(\sr_20_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[1]_net_1 ));
    DFN1E1C0 \sr_37_[9]  (.D(\sr_36_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[9]_net_1 ));
    DFN1E1C0 \sr_48_[10]  (.D(\sr_47_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[10]_net_1 ));
    DFN1E1C0 \sr_60_[5]  (.D(\sr_59_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[5]_net_1 ));
    DFN1E1C0 \sr_30_[5]  (.D(\sr_29_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[5]_net_1 ));
    DFN1E1C0 \sr_14_[4]  (.D(\sr_13_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[4]_net_1 ));
    DFN1E1C0 \sr_24_[8]  (.D(\sr_23_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[8]_net_1 ));
    DFN1E1C0 \sr_30_[4]  (.D(\sr_29_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[4]_net_1 ));
    DFN1E1C0 \sr_37_[6]  (.D(\sr_36_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[6]_net_1 ));
    DFN1E1C0 \sr_42_[6]  (.D(\sr_41_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[6]_net_1 ));
    DFN1E1C0 \sr_58_[4]  (.D(\sr_57_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[4]_net_1 ));
    DFN1E1C0 \sr_57_[10]  (.D(\sr_56_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[10]_net_1 ));
    DFN1E1C0 \sr_43_[7]  (.D(\sr_42_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[7]_net_1 ));
    DFN1E1C0 \sr_44_[2]  (.D(\sr_43_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[2]_net_1 ));
    DFN1E1C0 \sr_53_[7]  (.D(\sr_52_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[7]_net_1 ));
    DFN1E1C0 \sr_59_[1]  (.D(\sr_58_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[1]_net_1 ));
    DFN1E1C0 \sr_27_[10]  (.D(\sr_26_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[10]_net_1 ));
    DFN1E1C0 \sr_53_[8]  (.D(\sr_52_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[8]_net_1 ));
    DFN1E1C0 \sr_16_[4]  (.D(\sr_15_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[4]_net_1 ));
    DFN1E1C0 \sr_10_[11]  (.D(\sr_9_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[11]_net_1 ));
    DFN1E1C0 \sr_26_[8]  (.D(\sr_25_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[8]_net_1 ));
    DFN1E1C0 \sr_63_[7]  (.D(\sr_62_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[7]));
    DFN1E1C0 \sr_28_[7]  (.D(\sr_27_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[7]_net_1 ));
    DFN1E1C0 \sr_63_[8]  (.D(\sr_62_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[8]));
    DFN1E1C0 \sr_24_[0]  (.D(\sr_23_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[0]_net_1 ));
    DFN1E1C0 \sr_46_[2]  (.D(\sr_45_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[2]_net_1 ));
    DFN1E1C0 \sr_13_[5]  (.D(\sr_12_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[5]_net_1 ));
    DFN1E1C0 \sr_0_[2]  (.D(cur_error[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[2]));
    DFN1E1C0 \sr_0_[8]  (.D(cur_error[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[8]));
    DFN1E1C0 \sr_8_[3]  (.D(\sr_7_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[3]_net_1 ));
    DFN1E1C0 \sr_42_[11]  (.D(\sr_41_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[11]_net_1 ));
    DFN1E1C0 \sr_13_[3]  (.D(\sr_12_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[3]_net_1 ));
    DFN1E1C0 \sr_54_[10]  (.D(\sr_53_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[10]_net_1 ));
    DFN1E1C0 \sr_37_[11]  (.D(\sr_36_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[11]_net_1 ));
    DFN1E1C0 \sr_19_[7]  (.D(\sr_18_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[7]_net_1 ));
    DFN1E1C0 \sr_57_[1]  (.D(\sr_56_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[1]_net_1 ));
    DFN1E1C0 \sr_44_[11]  (.D(\sr_43_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[11]_net_1 ));
    DFN1E1C0 \sr_32_[10]  (.D(\sr_31_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[10]_net_1 ));
    DFN1E1C0 \sr_26_[0]  (.D(\sr_25_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[0]_net_1 ));
    DFN1E1C0 \sr_24_[10]  (.D(\sr_23_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[10]_net_1 ));
    DFN1E1C0 \sr_12_[1]  (.D(\sr_11_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[1]_net_1 ));
    DFN1E1C0 \sr_10_[4]  (.D(\sr_9_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[4]_net_1 ));
    DFN1E1C0 \sr_63_[0]  (.D(\sr_62_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[0]));
    DFN1E1C0 \sr_20_[8]  (.D(\sr_19_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[8]_net_1 ));
    DFN1E1C0 \sr_60_[12]  (.D(\sr_59_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[12]_net_1 ));
    DFN1E1C0 \sr_6_[10]  (.D(\sr_5_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[10]_net_1 ));
    DFN1E1C0 \sr_19_[6]  (.D(\sr_18_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[6]_net_1 ));
    DFN1E1C0 \sr_62_[5]  (.D(\sr_61_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[5]_net_1 ));
    DFN1E1C0 \sr_44_[8]  (.D(\sr_43_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[8]_net_1 ));
    DFN1E1C0 \sr_49_[5]  (.D(\sr_48_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[5]_net_1 ));
    DFN1E1C0 \sr_53_[0]  (.D(\sr_52_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[0]_net_1 ));
    DFN1E1C0 \sr_1_[2]  (.D(sr_new[2]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[2]));
    DFN1E1C0 \sr_40_[2]  (.D(\sr_39_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[2]_net_1 ));
    DFN1E1C0 \sr_32_[5]  (.D(\sr_31_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[5]_net_1 ));
    DFN1E1C0 \sr_1_[8]  (.D(sr_new[8]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[8]));
    DFN1E1C0 \sr_18_[12]  (.D(\sr_17_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[12]_net_1 ));
    DFN1E1C0 \sr_60_[10]  (.D(\sr_59_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[10]_net_1 ));
    DFN1E1C0 \sr_32_[4]  (.D(\sr_31_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[4]_net_1 ));
    DFN1E1C0 \sr_54_[3]  (.D(\sr_53_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[3]_net_1 ));
    DFN1E1C0 \sr_29_[9]  (.D(\sr_28_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[9]_net_1 ));
    DFN1E1C0 \sr_24_[2]  (.D(\sr_23_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[2]_net_1 ));
    DFN1E1C0 \sr_18_[9]  (.D(\sr_17_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[9]_net_1 ));
    DFN1E1C0 \sr_7_[9]  (.D(\sr_6_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[9]_net_1 ));
    DFN1E1C0 \sr_63_[10]  (.D(\sr_62_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[10]));
    DFN1E1C0 \sr_24_[5]  (.D(\sr_23_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[5]_net_1 ));
    DFN1E1C0 \sr_46_[8]  (.D(\sr_45_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[8]_net_1 ));
    DFN1E1C0 \sr_59_[11]  (.D(\sr_58_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[11]_net_1 ));
    DFN1E1C0 \sr_17_[7]  (.D(\sr_16_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[7]_net_1 ));
    DFN1E1C0 \sr_14_[8]  (.D(\sr_13_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[8]_net_1 ));
    DFN1E1C0 \sr_41_[3]  (.D(\sr_40_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[3]_net_1 ));
    DFN1E1C0 \sr_20_[0]  (.D(\sr_19_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[0]_net_1 ));
    DFN1E1C0 \sr_48_[0]  (.D(\sr_47_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[0]_net_1 ));
    DFN1E1C0 \sr_29_[1]  (.D(\sr_28_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[1]_net_1 ));
    DFN1E1C0 \sr_3_[10]  (.D(\sr_2_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[10]_net_1 ));
    DFN1E1C0 \sr_29_[11]  (.D(\sr_28_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[11]_net_1 ));
    DFN1E1C0 \sr_35_[1]  (.D(\sr_34_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[1]_net_1 ));
    DFN1E1C0 \sr_17_[6]  (.D(\sr_16_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[6]_net_1 ));
    DFN1E1C0 \sr_2_[3]  (.D(sr_prev[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[3]_net_1 ));
    DFN1E1C0 \sr_56_[3]  (.D(\sr_55_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[3]_net_1 ));
    DFN1E1C0 \sr_47_[5]  (.D(\sr_46_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[5]_net_1 ));
    DFN1E1C0 \sr_35_[2]  (.D(\sr_34_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[2]_net_1 ));
    DFN1E1C0 \sr_35_[12]  (.D(\sr_34_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[12]_net_1 ));
    DFN1E1C0 \sr_26_[2]  (.D(\sr_25_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[2]_net_1 ));
    DFN1E1C0 \sr_6_[2]  (.D(\sr_5_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[2]_net_1 ));
    DFN1E1C0 \sr_6_[8]  (.D(\sr_5_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[8]_net_1 ));
    DFN1E1C0 \sr_35_[7]  (.D(\sr_34_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[7]_net_1 ));
    DFN1E1C0 \sr_26_[5]  (.D(\sr_25_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[5]_net_1 ));
    DFN1E1C0 \sr_16_[8]  (.D(\sr_15_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[8]_net_1 ));
    DFN1E1C0 \sr_52_[12]  (.D(\sr_51_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[12]_net_1 ));
    DFN1E1C0 \sr_5_[2]  (.D(\sr_4_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[2]_net_1 ));
    DFN1E1C0 \sr_5_[8]  (.D(\sr_4_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[8]_net_1 ));
    DFN1E1C0 \sr_27_[9]  (.D(\sr_26_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[9]_net_1 ));
    DFN1E1C0 \sr_18_[11]  (.D(\sr_17_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[11]_net_1 ));
    DFN1E1C0 \sr_3_[9]  (.D(\sr_2_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[9]_net_1 ));
    DFN1E1C0 \sr_2_[11]  (.D(sr_prev[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[11]_net_1 ));
    DFN1E1C0 \sr_40_[8]  (.D(\sr_39_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[8]_net_1 ));
    DFN1E1C0 \sr_22_[12]  (.D(\sr_21_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[12]_net_1 ));
    DFN1E1C0 \sr_45_[9]  (.D(\sr_44_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[9]_net_1 ));
    DFN1E1C0 \sr_2_[12]  (.D(sr_prev[12]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[12]_net_1 ));
    DFN1E1C0 \sr_27_[1]  (.D(\sr_26_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[1]_net_1 ));
    DFN1E1C0 \sr_0__1[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_new_1_0));
    DFN1E1C0 \sr_9_[4]  (.D(\sr_8_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[4]_net_1 ));
    DFN1E1C0 \sr_12_[4]  (.D(\sr_11_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[4]_net_1 ));
    DFN1E1C0 \sr_56_[11]  (.D(\sr_55_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[11]_net_1 ));
    DFN1E1C0 \sr_22_[8]  (.D(\sr_21_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[8]_net_1 ));
    DFN1E1C0 \sr_14_[2]  (.D(\sr_13_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[2]_net_1 ));
    DFN1E1C0 \sr_46_[12]  (.D(\sr_45_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[12]_net_1 ));
    DFN1E1C0 \sr_50_[3]  (.D(\sr_49_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[3]_net_1 ));
    DFN1E1C0 \sr_20_[2]  (.D(\sr_19_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[2]_net_1 ));
    DFN1E1C0 \sr_44_[12]  (.D(\sr_43_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[12]_net_1 ));
    DFN1E1C0 \sr_26_[11]  (.D(\sr_25_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[11]_net_1 ));
    DFN1E1C0 \sr_14_[0]  (.D(\sr_13_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[0]_net_1 ));
    DFN1E1C0 \sr_34_[8]  (.D(\sr_33_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[8]_net_1 ));
    DFN1E1C0 \sr_20_[5]  (.D(\sr_19_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[5]_net_1 ));
    DFN1E1C0 \sr_10_[8]  (.D(\sr_9_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[8]_net_1 ));
    DFN1E1C0 \sr_42_[2]  (.D(\sr_41_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[2]_net_1 ));
    DFN1E1C0 \sr_55_[11]  (.D(\sr_54_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[11]_net_1 ));
    DFN1E1C0 \sr_51_[9]  (.D(\sr_50_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[9]_net_1 ));
    DFN1E1C0 \sr_54_[5]  (.D(\sr_53_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[5]_net_1 ));
    DFN1E1C0 \sr_25_[11]  (.D(\sr_24_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[11]_net_1 ));
    DFN1E1C0 \sr_21_[6]  (.D(\sr_20_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[6]_net_1 ));
    DFN1E1C0 \sr_57_[12]  (.D(\sr_56_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[12]_net_1 ));
    DFN1E1C0 \sr_16_[2]  (.D(\sr_15_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[2]_net_1 ));
    DFN1E1C0 \sr_35_[0]  (.D(\sr_34_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[0]_net_1 ));
    DFN1E1C0 \sr_16_[0]  (.D(\sr_15_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[0]_net_1 ));
    DFN1E1C0 \sr_36_[8]  (.D(\sr_35_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[8]_net_1 ));
    DFN1E1C0 \sr_27_[12]  (.D(\sr_26_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[12]_net_1 ));
    DFN1E1C0 \sr_22_[0]  (.D(\sr_21_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[0]_net_1 ));
    DFN1E1C0 \sr_0__0[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_new_0_0));
    DFN1E1C0 \sr_13_[11]  (.D(\sr_12_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[11]_net_1 ));
    DFN1E1C0 \sr_58_[10]  (.D(\sr_57_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[10]_net_1 ));
    DFN1E1C0 \sr_7_[12]  (.D(\sr_6_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[12]_net_1 ));
    DFN1E1C0 \sr_24_[3]  (.D(\sr_23_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[3]_net_1 ));
    DFN1E1C0 \sr_34_[9]  (.D(\sr_33_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[9]_net_1 ));
    DFN1E1C0 \sr_28_[10]  (.D(\sr_27_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[10]_net_1 ));
    DFN1E1C0 \sr_56_[5]  (.D(\sr_55_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[5]_net_1 ));
    DFN1E1C0 \sr_7_[10]  (.D(\sr_6_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[10]_net_1 ));
    DFN1E1C0 \sr_33_[1]  (.D(\sr_32_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[1]_net_1 ));
    DFN1E1C0 \sr_33_[2]  (.D(\sr_32_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[2]_net_1 ));
    DFN1E1C0 \sr_48_[7]  (.D(\sr_47_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[7]_net_1 ));
    DFN1E1C0 \sr_58_[7]  (.D(\sr_57_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[7]_net_1 ));
    DFN1E1C0 \sr_34_[6]  (.D(\sr_33_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[6]_net_1 ));
    DFN1E1C0 \sr_33_[7]  (.D(\sr_32_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[7]_net_1 ));
    DFN1E1C0 \sr_10_[2]  (.D(\sr_9_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[2]_net_1 ));
    DFN1E1C0 \sr_26_[3]  (.D(\sr_25_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[3]_net_1 ));
    DFN1E1C0 \sr_36_[9]  (.D(\sr_35_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[9]_net_1 ));
    DFN1E1C0 \sr_58_[8]  (.D(\sr_57_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[8]_net_1 ));
    DFN1E1C0 \sr_42_[8]  (.D(\sr_41_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[8]_net_1 ));
    DFN1E1C0 \sr_49_[3]  (.D(\sr_48_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[3]_net_1 ));
    DFN1E1C0 \sr_10_[0]  (.D(\sr_9_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[0]_net_1 ));
    DFN1E1C0 \sr_30_[8]  (.D(\sr_29_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[8]_net_1 ));
    DFN1E1C0 \sr_35_[10]  (.D(\sr_34_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[10]_net_1 ));
    DFN1E1C0 \sr_8_[4]  (.D(\sr_7_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[4]_net_1 ));
    DFN1E1C0 \sr_43_[12]  (.D(\sr_42_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[12]_net_1 ));
    DFN1E1C0 \sr_0_[9]  (.D(cur_error[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[9]));
    DFN1E1C0 \sr_43_[9]  (.D(\sr_42_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[9]_net_1 ));
    DFN1E1C0 \sr_50_[5]  (.D(\sr_49_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[5]_net_1 ));
    DFN1E1C0 \sr_52_[3]  (.D(\sr_51_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[3]_net_1 ));
    DFN1E1C0 \sr_22_[2]  (.D(\sr_21_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[2]_net_1 ));
    DFN1E1C0 \sr_18_[5]  (.D(\sr_17_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[5]_net_1 ));
    DFN1E1C0 \sr_7_[0]  (.D(\sr_6_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[0]_net_1 ));
    DFN1E1C0 \sr_36_[6]  (.D(\sr_35_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[6]_net_1 ));
    DFN1E1C0 \sr_60_[11]  (.D(\sr_59_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[11]_net_1 ));
    DFN1E1C0 \sr_45_[4]  (.D(\sr_44_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[4]_net_1 ));
    DFN1E1C0 \sr_22_[5]  (.D(\sr_21_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[5]_net_1 ));
    DFN1E1C0 \sr_35_[3]  (.D(\sr_34_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[3]_net_1 ));
    DFN1E1C0 \sr_7_[6]  (.D(\sr_6_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[6]_net_1 ));
    DFN1E1C0 \sr_12_[8]  (.D(\sr_11_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[8]_net_1 ));
    DFN1E1C0 \sr_55_[6]  (.D(\sr_54_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[6]_net_1 ));
    DFN1E1C0 \sr_52_[11]  (.D(\sr_51_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[11]_net_1 ));
    DFN1E1C0 \sr_18_[3]  (.D(\sr_17_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[3]_net_1 ));
    DFN1E1C0 \sr_36_[10]  (.D(\sr_35_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[10]_net_1 ));
    DFN1E1C0 \sr_25_[4]  (.D(\sr_24_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[4]_net_1 ));
    DFN1E1C0 \sr_22_[11]  (.D(\sr_21_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[11]_net_1 ));
    DFN1E1C0 \sr_20_[3]  (.D(\sr_19_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[3]_net_1 ));
    DFN1E1C0 \sr_30_[9]  (.D(\sr_29_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[9]_net_1 ));
    DFN1E1C0 \sr_47_[3]  (.D(\sr_46_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[3]_net_1 ));
    DFN1E1C0 \sr_54_[11]  (.D(\sr_53_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[11]_net_1 ));
    DFN1E1C0 \sr_4_[7]  (.D(\sr_3_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[7]_net_1 ));
    DFN1E1C0 \sr_31_[12]  (.D(\sr_30_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[12]_net_1 ));
    DFN1E1C0 \sr_54_[1]  (.D(\sr_53_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[1]_net_1 ));
    DFN1E1C0 \sr_24_[11]  (.D(\sr_23_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[11]_net_1 ));
    DFN1E1C0 \sr_1_[9]  (.D(sr_new[9]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[9]));
    DFN1E1C0 \sr_58_[0]  (.D(\sr_57_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[0]_net_1 ));
    DFN1E1C0 \sr_33_[0]  (.D(\sr_32_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[0]_net_1 ));
    DFN1E1C0 \sr_41_[1]  (.D(\sr_40_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[1]_net_1 ));
    DFN1E1C0 \sr_30_[6]  (.D(\sr_29_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[6]_net_1 ));
    DFN1E1C0 \sr_7_[1]  (.D(\sr_6_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[1]_net_1 ));
    DFN1E1C0 \sr_3_[0]  (.D(\sr_2_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[0]_net_1 ));
    DFN1E1C0 \sr_45_[6]  (.D(\sr_44_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[6]_net_1 ));
    DFN1E1C0 \sr_3_[6]  (.D(\sr_2_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[6]_net_1 ));
    DFN1E1C0 \sr_59_[9]  (.D(\sr_58_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[9]_net_1 ));
    DFN1E1C0 \sr_2_[4]  (.D(sr_prev[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[4]_net_1 ));
    DFN1E1C0 \sr_56_[1]  (.D(\sr_55_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[1]_net_1 ));
    DFN1E1C0 \sr_29_[6]  (.D(\sr_28_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[6]_net_1 ));
    DFN1E1C0 \sr_9_[2]  (.D(\sr_8_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[2]_net_1 ));
    DFN1E1C0 \sr_9_[8]  (.D(\sr_8_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[8]_net_1 ));
    DFN1E1C0 \sr_17_[11]  (.D(\sr_16_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[11]_net_1 ));
    DFN1E1C0 \sr_12_[2]  (.D(\sr_11_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[2]_net_1 ));
    DFN1E1C0 \sr_12_[10]  (.D(\sr_11_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[10]_net_1 ));
    DFN1E1C0 \sr_12_[0]  (.D(\sr_11_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[0]_net_1 ));
    DFN1E1C0 \sr_32_[8]  (.D(\sr_31_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[8]_net_1 ));
    DFN1E1C0 \sr_14_[7]  (.D(\sr_13_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[7]_net_1 ));
    DFN1E1C0 \sr_6_[9]  (.D(\sr_5_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[9]_net_1 ));
    DFN1E1C0 \sr_31_[10]  (.D(\sr_30_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[10]_net_1 ));
    DFN1E1C0 \sr_31_[11]  (.D(\sr_30_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[11]_net_1 ));
    DFN1E1C0 \sr_14_[6]  (.D(\sr_13_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[6]_net_1 ));
    DFN1E1C0 \sr_5_[10]  (.D(\sr_4_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[10]_net_1 ));
    DFN1E1C0 \sr_5_[9]  (.D(\sr_4_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[9]_net_1 ));
    DFN1E1C0 \sr_52_[5]  (.D(\sr_51_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[5]_net_1 ));
    DFN1E1C0 \sr_3_[1]  (.D(\sr_2_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[1]_net_1 ));
    DFN1E1C0 \sr_44_[5]  (.D(\sr_43_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[5]_net_1 ));
    DFN1E1C0 \sr_57_[9]  (.D(\sr_56_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[9]_net_1 ));
    DFN1E1C0 \sr_50_[1]  (.D(\sr_49_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[1]_net_1 ));
    DFN1E1C0 \sr_16_[7]  (.D(\sr_15_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[7]_net_1 ));
    DFN1E1C0 \sr_51_[2]  (.D(\sr_50_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[2]_net_1 ));
    DFN1E1C0 \sr_27_[6]  (.D(\sr_26_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[6]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1C0 \sr_43_[4]  (.D(\sr_42_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[4]_net_1 ));
    DFN1E1C0 \sr_24_[9]  (.D(\sr_23_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[9]_net_1 ));
    DFN1E1C0 \sr_22_[3]  (.D(\sr_21_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[3]_net_1 ));
    DFN1E1C0 \sr_33_[3]  (.D(\sr_32_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[3]_net_1 ));
    DFN1E1C0 \sr_32_[9]  (.D(\sr_31_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[9]_net_1 ));
    DFN1E1C0 \sr_15_[1]  (.D(\sr_14_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[1]_net_1 ));
    DFN1E1C0 \sr_53_[6]  (.D(\sr_52_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[6]_net_1 ));
    DFN1E1C0 \sr_60_[1]  (.D(\sr_59_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[1]_net_1 ));
    DFN1E1C0 \sr_16_[6]  (.D(\sr_15_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[6]_net_1 ));
    DFN1E1C0 \sr_61_[2]  (.D(\sr_60_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[2]_net_1 ));
    DFN1E1C0 \sr_23_[4]  (.D(\sr_22_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[4]_net_1 ));
    DFN1E1C0 \sr_46_[5]  (.D(\sr_45_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[5]_net_1 ));
    DFN1E1C0 \sr_24_[1]  (.D(\sr_23_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[1]_net_1 ));
    DFN1E1C0 \sr_63_[6]  (.D(\sr_62_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[6]));
    DFN1E1C0 \sr_49_[12]  (.D(\sr_48_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[12]_net_1 ));
    DFN1E1C0 \sr_56_[12]  (.D(\sr_55_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[12]_net_1 ));
    DFN1E1C0 \sr_54_[12]  (.D(\sr_53_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[12]_net_1 ));
    DFN1E1C0 \sr_35_[5]  (.D(\sr_34_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[5]_net_1 ));
    DFN1E1C0 \sr_15_[12]  (.D(\sr_14_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[12]_net_1 ));
    DFN1E1C0 \sr_32_[6]  (.D(\sr_31_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[6]_net_1 ));
    DFN1E1C0 \sr_26_[12]  (.D(\sr_25_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[12]_net_1 ));
    DFN1E1C0 \sr_35_[4]  (.D(\sr_34_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[4]_net_1 ));
    DFN1E1C0 \sr_26_[9]  (.D(\sr_25_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[9]_net_1 ));
    DFN1E1C0 \sr_24_[12]  (.D(\sr_23_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[12]_net_1 ));
    DFN1E1C0 \sr_51_[4]  (.D(\sr_50_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[4]_net_1 ));
    DFN1E1C0 \sr_10_[7]  (.D(\sr_9_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[7]_net_1 ));
    DFN1E1C0 \sr_8_[2]  (.D(\sr_7_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[2]_net_1 ));
    DFN1E1C0 \sr_40_[12]  (.D(\sr_39_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[12]_net_1 ));
    DFN1E1C0 \sr_8_[8]  (.D(\sr_7_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[8]_net_1 ));
    DFN1E1C0 \sr_26_[1]  (.D(\sr_25_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[1]_net_1 ));
    DFN1E1C0 \sr_61_[4]  (.D(\sr_60_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[4]_net_1 ));
    DFN1E1C0 \sr_0_[0]  (.D(cur_error[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[0]));
    DFN1E1C0 \sr_43_[6]  (.D(\sr_42_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[6]_net_1 ));
    DFN1E1C0 \sr_10_[6]  (.D(\sr_9_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[6]_net_1 ));
    DFN1E1C0 \sr_21_[7]  (.D(\sr_20_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[7]_net_1 ));
    DFN1E1C0 \sr_0_[6]  (.D(cur_error[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[6]));
    DFN1E1C0 \sr_40_[5]  (.D(\sr_39_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[5]_net_1 ));
    DFN1E1C0 \sr_40_[10]  (.D(\sr_39_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[10]_net_1 ));
    DFN1E1C0 \sr_43_[10]  (.D(\sr_42_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[10]_net_1 ));
    DFN1E1C0 \sr_38_[1]  (.D(\sr_37_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[1]_net_1 ));
    DFN1E1C0 \sr_49_[1]  (.D(\sr_48_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[1]_net_1 ));
    DFN1E1C0 \sr_63_[11]  (.D(\sr_62_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[11]));
    DFN1E1C0 \sr_20_[9]  (.D(\sr_19_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[9]_net_1 ));
    DFN1E1C0 \sr_38_[2]  (.D(\sr_37_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[2]_net_1 ));
    DFN1E1C0 \sr_38_[7]  (.D(\sr_37_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[7]_net_1 ));
    DFN1E1C0 \sr_52_[1]  (.D(\sr_51_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[1]_net_1 ));
    DFN1E1C0 \sr_20_[1]  (.D(\sr_19_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[1]_net_1 ));
    DFN1E1C0 \sr_1_[0]  (.D(sr_new[0]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[0]));
    DFN1E1C0 \sr_61_[9]  (.D(\sr_60_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[9]_net_1 ));
    DFN1E1C0 \sr_0_[1]  (.D(cur_error[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[1]));
    DFN1E1C0 \sr_15_[4]  (.D(\sr_14_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[4]_net_1 ));
    DFN1E1C0 \sr_1_[6]  (.D(sr_new[6]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[6]));
    DFN1E1C0 \sr_62_[1]  (.D(\sr_61_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[1]_net_1 ));
    DFN1E1C0 \sr_25_[8]  (.D(\sr_24_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[8]_net_1 ));
    DFN1E1C0 \sr_48_[9]  (.D(\sr_47_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[9]_net_1 ));
    DFN1E1C0 \sr_1_[11]  (.D(sr_new[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_prev[11]));
    DFN1E1C0 \sr_49_[10]  (.D(\sr_48_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[10]_net_1 ));
    DFN1E1C0 \sr_53_[12]  (.D(\sr_52_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[12]_net_1 ));
    DFN1E1C0 \sr_13_[1]  (.D(\sr_12_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[1]_net_1 ));
    DFN1E1C0 \sr_7_[5]  (.D(\sr_6_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[5]_net_1 ));
    DFN1E1C0 \sr_5_[12]  (.D(\sr_4_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[12]_net_1 ));
    DFN1E1C0 \sr_47_[1]  (.D(\sr_46_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[1]_net_1 ));
    DFN1E1C0 \sr_23_[12]  (.D(\sr_22_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[12]_net_1 ));
    DFN1E1C0 \sr_63_[5]  (.D(\sr_62_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[5]));
    DFN1E1C0 \sr_45_[2]  (.D(\sr_44_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[2]_net_1 ));
    DFN1E1C0 \sr_2_[2]  (.D(sr_prev[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[2]_net_1 ));
    DFN1E1C0 \sr_2_[8]  (.D(sr_prev[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[8]_net_1 ));
    DFN1E1C0 \sr_11_[9]  (.D(\sr_10_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[9]_net_1 ));
    DFN1E1C0 \sr_33_[5]  (.D(\sr_32_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[5]_net_1 ));
    DFN1E1C0 \sr_59_[2]  (.D(\sr_58_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[2]_net_1 ));
    DFN1E1C0 \sr_12_[7]  (.D(\sr_11_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[7]_net_1 ));
    DFN1E1C0 \sr_6_[0]  (.D(\sr_5_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[0]_net_1 ));
    DFN1E1C0 \sr_41_[0]  (.D(\sr_40_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[0]_net_1 ));
    DFN1E1C0 \sr_1_[1]  (.D(sr_new[1]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[1]));
    DFN1E1C0 \sr_33_[4]  (.D(\sr_32_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[4]_net_1 ));
    DFN1E1C0 \sr_9_[12]  (.D(\sr_8_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[12]_net_1 ));
    DFN1E1C0 \sr_25_[0]  (.D(\sr_24_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[0]_net_1 ));
    DFN1E1C0 \sr_6_[6]  (.D(\sr_5_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[6]_net_1 ));
    DFN1E1C0 \sr_15_[10]  (.D(\sr_14_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[10]_net_1 ));
    DFN1E1C0 \sr_12_[6]  (.D(\sr_11_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[6]_net_1 ));
    DFN1E1C0 \sr_61_[3]  (.D(\sr_60_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[3]_net_1 ));
    DFN1E1C0 \sr_5_[0]  (.D(\sr_4_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[0]_net_1 ));
    DFN1E1C0 \sr_44_[3]  (.D(\sr_43_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[3]_net_1 ));
    DFN1E1C0 \sr_38_[0]  (.D(\sr_37_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[0]_net_1 ));
    DFN1E1C0 \sr_42_[5]  (.D(\sr_41_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[5]_net_1 ));
    DFN1E1C0 \sr_5_[6]  (.D(\sr_4_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[6]_net_1 ));
    DFN1E1C0 \sr_3_[5]  (.D(\sr_2_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[5]_net_1 ));
    DFN1E1C0 \sr_4_[3]  (.D(\sr_3_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[3]_net_1 ));
    DFN1E1C0 \sr_9_[9]  (.D(\sr_8_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[9]_net_1 ));
    DFN1E1C0 \sr_37_[10]  (.D(\sr_36_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[10]_net_1 ));
    DFN1E1C0 \sr_22_[9]  (.D(\sr_21_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[9]_net_1 ));
    DFN1E1C0 \sr_59_[4]  (.D(\sr_58_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[4]_net_1 ));
    DFN1E1C0 \sr_16_[10]  (.D(\sr_15_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[10]_net_1 ));
    DFN1E1C0 \sr_57_[2]  (.D(\sr_56_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[2]_net_1 ));
    DFN1E1C0 \sr_46_[3]  (.D(\sr_45_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[3]_net_1 ));
    DFN1E1C0 \sr_6_[1]  (.D(\sr_5_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[1]_net_1 ));
    DFN1E1C0 \sr_45_[8]  (.D(\sr_44_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[8]_net_1 ));
    DFN1E1C0 \sr_22_[1]  (.D(\sr_21_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[1]_net_1 ));
    DFN1E1C0 \sr_29_[7]  (.D(\sr_28_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[7]_net_1 ));
    DFN1E1C0 \sr_11_[12]  (.D(\sr_10_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[12]_net_1 ));
    DFN1E1C0 \sr_5_[1]  (.D(\sr_4_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[1]_net_1 ));
    DFN1E1C0 \sr_4_[10]  (.D(\sr_3_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[10]_net_1 ));
    DFN1E1C0 \sr_55_[3]  (.D(\sr_54_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[3]_net_1 ));
    DFN1E1C0 \sr_25_[2]  (.D(\sr_24_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[2]_net_1 ));
    DFN1E1C0 \sr_13_[4]  (.D(\sr_12_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[4]_net_1 ));
    DFN1E1C0 \sr_62_[10]  (.D(\sr_61_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[10]_net_1 ));
    DFN1E1C0 \sr_23_[8]  (.D(\sr_22_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[8]_net_1 ));
    DFN1E1C0 \sr_25_[5]  (.D(\sr_24_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[5]_net_1 ));
    DFN1E1C0 \sr_15_[8]  (.D(\sr_14_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[8]_net_1 ));
    DFN1E1C0 \sr_34_[10]  (.D(\sr_33_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[10]_net_1 ));
    DFN1E1C0 \sr_57_[4]  (.D(\sr_56_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[4]_net_1 ));
    DFN1E1C0 \sr_40_[3]  (.D(\sr_39_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[3]_net_1 ));
    DFN1E1C0 \sr_48_[4]  (.D(\sr_47_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[4]_net_1 ));
    DFN1E1C0 \sr_38_[3]  (.D(\sr_37_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[3]_net_1 ));
    DFN1E1C0 \sr_43_[2]  (.D(\sr_42_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[2]_net_1 ));
    DFN1E1C0 \sr_58_[6]  (.D(\sr_57_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[6]_net_1 ));
    DFN1E1C0 \sr_54_[9]  (.D(\sr_53_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[9]_net_1 ));
    DFN1E1C0 \sr_28_[4]  (.D(\sr_27_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[4]_net_1 ));
    DFN1E1C0 \sr_27_[7]  (.D(\sr_26_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[7]_net_1 ));
    DFN1E1C0 \sr_24_[6]  (.D(\sr_23_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[6]_net_1 ));
    DFN1E1C0 \sr_40_[11]  (.D(\sr_39_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[11]_net_1 ));
    DFN1E1C0 \sr_11_[10]  (.D(\sr_10_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[10]_net_1 ));
    DFN1E1C0 \sr_23_[0]  (.D(\sr_22_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[0]_net_1 ));
    DFN1E1C0 \sr_11_[11]  (.D(\sr_10_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[11]_net_1 ));
    DFN1E1C0 \sr_59_[12]  (.D(\sr_58_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[12]_net_1 ));
    DFN1E1C0 \sr_8_[9]  (.D(\sr_7_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[9]_net_1 ));
    DFN1E1C0 \sr_1_[10]  (.D(sr_new[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_prev[10]));
    DFN1E1C0 \sr_41_[7]  (.D(\sr_40_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[7]_net_1 ));
    DFN1E1C0 \sr_29_[12]  (.D(\sr_28_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[12]_net_1 ));
    DFN1E1C0 \sr_19_[9]  (.D(\sr_18_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[9]_net_1 ));
    DFN1E1C0 \sr_56_[9]  (.D(\sr_55_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[9]_net_1 ));
    DFN1E1C0 \sr_51_[7]  (.D(\sr_50_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[7]_net_1 ));
    DFN1E1C0 \sr_39_[11]  (.D(\sr_38_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[11]_net_1 ));
    DFN1E1C0 \sr_26_[6]  (.D(\sr_25_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[6]_net_1 ));
    DFN1E1C0 \sr_51_[8]  (.D(\sr_50_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[8]_net_1 ));
    DFN1E1C0 \sr_50_[12]  (.D(\sr_49_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[12]_net_1 ));
    DFN1E1C0 \sr_49_[0]  (.D(\sr_48_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[0]_net_1 ));
    DFN1E1C0 \sr_0_[5]  (.D(cur_error[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[5]));
    DFN1E1C0 \sr_15_[2]  (.D(\sr_14_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[2]_net_1 ));
    DFN1E1C0 \sr_61_[7]  (.D(\sr_60_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[7]_net_1 ));
    DFN1E1C0 \sr_48_[6]  (.D(\sr_47_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[6]_net_1 ));
    DFN1E1C0 \sr_15_[0]  (.D(\sr_14_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[0]_net_1 ));
    DFN1E1C0 \sr_35_[8]  (.D(\sr_34_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[8]_net_1 ));
    DFN1E1C0 \sr_61_[8]  (.D(\sr_60_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[8]_net_1 ));
    DFN1E1C0 \sr_20_[12]  (.D(\sr_19_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[12]_net_1 ));
    DFN1E1C0 \sr_43_[8]  (.D(\sr_42_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[8]_net_1 ));
    DFN1E1C0 \sr_11_[5]  (.D(\sr_10_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[5]_net_1 ));
    DFN1E1C0 \sr_50_[10]  (.D(\sr_49_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[10]_net_1 ));
    DFN1E1C0 \sr_55_[5]  (.D(\sr_54_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[5]_net_1 ));
    DFN1E1C0 \sr_53_[10]  (.D(\sr_52_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[10]_net_1 ));
    DFN1E1C0 \sr_48_[12]  (.D(\sr_47_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[12]_net_1 ));
    DFN1E1C0 \sr_32_[12]  (.D(\sr_31_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[12]_net_1 ));
    DFN1E1C0 \sr_11_[3]  (.D(\sr_10_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[3]_net_1 ));
    DFN1E1C0 \sr_0_[11]  (.D(cur_error[11]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable), .Q(sr_new[11]));
    DFN1E1C0 \sr_20_[10]  (.D(\sr_19_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[10]_net_1 ));
    DFN1E1C0 \sr_50_[9]  (.D(\sr_49_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[9]_net_1 ));
    DFN1E1C0 \sr_17_[9]  (.D(\sr_16_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[9]_net_1 ));
    DFN1E1C0 \sr_23_[10]  (.D(\sr_22_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[10]_net_1 ));
    DFN1E1C0 \sr_20_[6]  (.D(\sr_19_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[6]_net_1 ));
    DFN1E1C0 \sr_53_[3]  (.D(\sr_52_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[3]_net_1 ));
    DFN1E1C0 \sr_23_[2]  (.D(\sr_22_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[2]_net_1 ));
    DFN1E1C0 \sr_1_[5]  (.D(sr_new[5]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[5]));
    DFN1E1C0 \sr_61_[0]  (.D(\sr_60_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[0]_net_1 ));
    DFN1E1C0 \sr_47_[0]  (.D(\sr_46_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[0]_net_1 ));
    DFN1E1C0 \sr_23_[5]  (.D(\sr_22_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[5]_net_1 ));
    DFN1E1C0 \sr_42_[3]  (.D(\sr_41_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[3]_net_1 ));
    DFN1E1C0 \sr_25_[3]  (.D(\sr_24_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[3]_net_1 ));
    DFN1E1C0 \sr_35_[9]  (.D(\sr_34_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[9]_net_1 ));
    DFN1E1C0 \sr_13_[8]  (.D(\sr_12_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[8]_net_1 ));
    DFN1E1C0 \sr_36_[11]  (.D(\sr_35_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[11]_net_1 ));
    DFN1E1C0 \sr_51_[0]  (.D(\sr_50_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[0]_net_1 ));
    DFN1E1C0 \sr_18_[1]  (.D(\sr_17_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[1]_net_1 ));
    DFN1E1C0 \sr_2_[9]  (.D(sr_prev[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[9]_net_1 ));
    DFN1E1C0 \sr_9_[0]  (.D(\sr_8_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[0]_net_1 ));
    DFN1E1C0 \sr_59_[10]  (.D(\sr_58_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[10]_net_1 ));
    DFN1E1C0 \sr_35_[11]  (.D(\sr_34_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[11]_net_1 ));
    DFN1E1C0 \sr_35_[6]  (.D(\sr_34_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[6]_net_1 ));
    DFN1E1C0 \sr_9_[6]  (.D(\sr_8_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[6]_net_1 ));
    DFN1E1C0 \sr_29_[10]  (.D(\sr_28_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[10]_net_1 ));
    DFN1E1C0 \sr_44_[1]  (.D(\sr_43_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[1]_net_1 ));
    DFN1E1C0 \sr_38_[5]  (.D(\sr_37_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[5]_net_1 ));
    DFN1E1C0 \sr_37_[12]  (.D(\sr_36_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[12]_net_1 ));
    DFN1E1C0 \sr_6_[5]  (.D(\sr_5_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[5]_net_1 ));
    DFN1E1C0 \sr_48_[11]  (.D(\sr_47_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[11]_net_1 ));
    DFN1E1C0 \sr_38_[4]  (.D(\sr_37_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[4]_net_1 ));
    DFN1E1C0 \sr_4_[4]  (.D(\sr_3_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[4]_net_1 ));
    DFN1E1C0 \sr_38_[10]  (.D(\sr_37_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[10]_net_1 ));
    DFN1E1C0 \sr_5_[5]  (.D(\sr_4_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[5]_net_1 ));
    DFN1E1C0 \sr_13_[2]  (.D(\sr_12_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[2]_net_1 ));
    DFN1E1C0 \sr_46_[1]  (.D(\sr_45_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[1]_net_1 ));
    DFN1E1C0 \sr_9_[1]  (.D(\sr_8_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[1]_net_1 ));
    DFN1E1C0 \sr_13_[0]  (.D(\sr_12_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[0]_net_1 ));
    DFN1E1C0 \sr_33_[8]  (.D(\sr_32_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[8]_net_1 ));
    DFN1E1C0 \sr_49_[7]  (.D(\sr_48_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[7]_net_1 ));
    DFN1E1C0 \sr_59_[7]  (.D(\sr_58_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[7]_net_1 ));
    DFN1E1C0 \sr_52_[9]  (.D(\sr_51_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[9]_net_1 ));
    DFN1E1C0 \sr_59_[8]  (.D(\sr_58_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[8]_net_1 ));
    DFN1E1C0 \sr_53_[5]  (.D(\sr_52_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[5]_net_1 ));
    DFN1E1C0 \sr_22_[6]  (.D(\sr_21_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[6]_net_1 ));
    DFN1E1C0 \sr_55_[1]  (.D(\sr_54_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[1]_net_1 ));
    DFN1E1C0 \sr_54_[2]  (.D(\sr_53_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[2]_net_1 ));
    DFN1E1C0 \sr_43_[11]  (.D(\sr_42_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[11]_net_1 ));
    DFN1E1C0 \sr_8_[0]  (.D(\sr_7_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[0]_net_1 ));
    DFN1E1C0 \sr_23_[3]  (.D(\sr_22_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[3]_net_1 ));
    DFN1E1C0 \sr_40_[1]  (.D(\sr_39_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[1]_net_1 ));
    DFN1E1C0 \sr_33_[9]  (.D(\sr_32_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[9]_net_1 ));
    DFN1E1C0 \sr_19_[5]  (.D(\sr_18_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[5]_net_1 ));
    DFN1E1C0 \sr_18_[4]  (.D(\sr_17_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[4]_net_1 ));
    DFN1E1C0 \sr_28_[8]  (.D(\sr_27_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[8]_net_1 ));
    DFN1E1C0 \sr_8_[6]  (.D(\sr_7_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[6]_net_1 ));
    DFN1E1C0 \sr_32_[11]  (.D(\sr_31_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[11]_net_1 ));
    DFN1E1C0 \sr_61_[12]  (.D(\sr_60_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[12]_net_1 ));
    DFN1E1C0 \sr_19_[3]  (.D(\sr_18_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[3]_net_1 ));
    DFN1E1C0 \sr_8_[11]  (.D(\sr_7_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[11]_net_1 ));
    DFN1E1C0 \sr_47_[7]  (.D(\sr_46_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[7]_net_1 ));
    DFN1E1C0 \sr_57_[7]  (.D(\sr_56_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[7]_net_1 ));
    DFN1E1C0 \sr_56_[2]  (.D(\sr_55_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[2]_net_1 ));
    DFN1E1C0 \sr_17_[10]  (.D(\sr_16_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[10]_net_1 ));
    DFN1E1C0 \sr_57_[8]  (.D(\sr_56_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[8]_net_1 ));
    DFN1E1C0 \sr_48_[2]  (.D(\sr_47_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[2]_net_1 ));
    DFN1E1C0 \sr_15_[7]  (.D(\sr_14_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[7]_net_1 ));
    DFN1E1C0 \sr_34_[11]  (.D(\sr_33_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[11]_net_1 ));
    DFN1E1C0 \sr_33_[6]  (.D(\sr_32_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[6]_net_1 ));
    DFN1E1C0 \sr_54_[4]  (.D(\sr_53_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[4]_net_1 ));
    DFN1E1C0 \sr_15_[6]  (.D(\sr_14_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[6]_net_1 ));
    DFN1E1C0 \sr_59_[0]  (.D(\sr_58_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[0]_net_1 ));
    DFN1E1C0 \sr_50_[11]  (.D(\sr_49_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[11]_net_1 ));
    DFN1E1C0 \sr_45_[5]  (.D(\sr_44_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[5]_net_1 ));
    DFN1E1C0 \sr_8_[1]  (.D(\sr_7_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[1]_net_1 ));
    DFN1E1C0 \sr_31_[1]  (.D(\sr_30_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[1]_net_1 ));
    DFN1E1C0 \sr_28_[0]  (.D(\sr_27_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[0]_net_1 ));
    DFN1E1C0 \sr_17_[5]  (.D(\sr_16_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[5]_net_1 ));
    DFN1E1C0 \sr_24_[7]  (.D(\sr_23_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[7]_net_1 ));
    DFN1E1C0 \sr_20_[11]  (.D(\sr_19_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[11]_net_1 ));
    DFN1E1C0 \sr_31_[2]  (.D(\sr_30_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[2]_net_1 ));
    DFN1E1C0 \sr_17_[3]  (.D(\sr_16_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[3]_net_1 ));
    DFN1E1C0 \sr_56_[4]  (.D(\sr_55_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[4]_net_1 ));
    DFN1E1C0 \sr_31_[7]  (.D(\sr_30_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[7]_net_1 ));
    DFN1E1C0 \sr_25_[9]  (.D(\sr_24_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[9]_net_1 ));
    DFN1E1C0 \sr_61_[10]  (.D(\sr_60_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[10]_net_1 ));
    DFN1E1C0 \sr_50_[2]  (.D(\sr_49_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[2]_net_1 ));
    DFN1E1C0 \sr_14_[10]  (.D(\sr_13_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[10]_net_1 ));
    DFN1E1C0 \sr_61_[11]  (.D(\sr_60_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[11]_net_1 ));
    DFN1E1C0 \sr_25_[1]  (.D(\sr_24_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[1]_net_1 ));
    DFN1E1C0 \sr_60_[2]  (.D(\sr_59_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[2]_net_1 ));
    DFN1E1C0 \sr_26_[7]  (.D(\sr_25_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[7]_net_1 ));
    DFN1E1C0 \sr_2_[0]  (.D(sr_prev[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[0]_net_1 ));
    DFN1E1C0 \sr_41_[9]  (.D(\sr_40_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[9]_net_1 ));
    DFN1E1C0 \sr_57_[0]  (.D(\sr_56_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[0]_net_1 ));
    DFN1E1C0 \sr_48_[8]  (.D(\sr_47_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[8]_net_1 ));
    DFN1E1C0 \sr_53_[1]  (.D(\sr_52_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[1]_net_1 ));
    DFN1E1C0 \sr_2_[6]  (.D(sr_prev[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[6]_net_1 ));
    DFN1E1C0 \sr_7_[7]  (.D(\sr_6_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[7]_net_1 ));
    DFN1E1C0 \sr_42_[1]  (.D(\sr_41_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[1]_net_1 ));
    DFN1E1C0 \sr_63_[1]  (.D(\sr_62_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[1]));
    DFN1E1C0 \sr_50_[4]  (.D(\sr_49_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[4]_net_1 ));
    DFN1E1C0 \sr_58_[12]  (.D(\sr_57_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[12]_net_1 ));
    DFN1E1C0 \sr_58_[3]  (.D(\sr_57_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[3]_net_1 ));
    DFN1E1C0 \sr_28_[2]  (.D(\sr_27_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[2]_net_1 ));
    DFN1E1C0 \sr_4_[2]  (.D(\sr_3_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[2]_net_1 ));
    DFN1E1C0 \sr_4_[8]  (.D(\sr_3_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[8]_net_1 ));
    DFN1E1C0 \sr_28_[5]  (.D(\sr_27_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[5]_net_1 ));
    DFN1E1C0 \sr_28_[12]  (.D(\sr_27_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[12]_net_1 ));
    DFN1E1C0 \sr_60_[4]  (.D(\sr_59_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[4]_net_1 ));
    DFN1E1C0 \sr_19_[11]  (.D(\sr_18_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[11]_net_1 ));
    DFN1E1C0 \sr_14_[9]  (.D(\sr_13_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[9]_net_1 ));
    DFN1E1C0 \sr_18_[8]  (.D(\sr_17_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[8]_net_1 ));
    DFN1E1C0 \sr_47_[11]  (.D(\sr_46_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[11]_net_1 ));
    DFN1E1C0 \sr_20_[7]  (.D(\sr_19_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[7]_net_1 ));
    DFN1E1C0 \sr_2_[1]  (.D(sr_prev[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[1]_net_1 ));
    DFN1E1C0 \sr_31_[0]  (.D(\sr_30_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[0]_net_1 ));
    DFN1E1C0 \sr_42_[10]  (.D(\sr_41_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[10]_net_1 ));
    DFN1E1C0 \sr_44_[0]  (.D(\sr_43_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[0]_net_1 ));
    DFN1E1C0 \sr_13_[7]  (.D(\sr_12_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[7]_net_1 ));
    DFN1E1C0 \sr_36_[12]  (.D(\sr_35_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[12]_net_1 ));
    DFN1E1C0 \sr_9_[5]  (.D(\sr_8_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[5]_net_1 ));
    DFN1E1C0 \sr_34_[12]  (.D(\sr_33_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[12]_net_1 ));
    DFN1E1C0 \sr_3_[7]  (.D(\sr_2_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[7]_net_1 ));
    DFN1E1C0 \sr_13_[6]  (.D(\sr_12_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[6]_net_1 ));
    DFN1E1C0 \sr_16_[9]  (.D(\sr_15_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[9]_net_1 ));
    DFN1E1C0 \sr_12_[12]  (.D(\sr_11_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[12]_net_1 ));
    DFN1E1C0 \sr_43_[5]  (.D(\sr_42_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[5]_net_1 ));
    DFN1E1C0 \sr_46_[0]  (.D(\sr_45_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[0]_net_1 ));
    DFN1E1C0 \sr_52_[2]  (.D(\sr_51_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[2]_net_1 ));
    DFN1E1C0 \sr_60_[9]  (.D(\sr_59_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[9]_net_1 ));
    DFN1E1C0 \sr_4_[12]  (.D(\sr_3_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[12]_net_1 ));
    DFN1E1C0 \sr_58_[11]  (.D(\sr_57_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[11]_net_1 ));
    DFN1E1C0 \sr_3_[12]  (.D(\sr_2_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[12]_net_1 ));
    DFN1E1C0 \sr_23_[9]  (.D(\sr_22_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[9]_net_1 ));
    DFN1E1C0 \sr_28_[11]  (.D(\sr_27_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[11]_net_1 ));
    DFN1E1C0 \sr_62_[2]  (.D(\sr_61_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[2]_net_1 ));
    DFN1E1C0 \sr_16_[11]  (.D(\sr_15_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[11]_net_1 ));
    DFN1E1C0 \sr_1_[12]  (.D(sr_new_0_0), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_prev[12]));
    DFN1E1C0 \sr_18_[2]  (.D(\sr_17_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[2]_net_1 ));
    DFN1E1C0 \sr_39_[1]  (.D(\sr_38_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[1]_net_1 ));
    DFN1E1C0 \sr_23_[1]  (.D(\sr_22_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[1]_net_1 ));
    DFN1E1C0 \sr_18_[0]  (.D(\sr_17_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[0]_net_1 ));
    DFN1E1C0 \sr_38_[8]  (.D(\sr_37_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[8]_net_1 ));
    DFN1E1C0 \sr_8_[10]  (.D(\sr_7_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[10]_net_1 ));
    DFN1E1C0 \sr_10_[9]  (.D(\sr_9_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[9]_net_1 ));
    DFN1E1C0 \sr_45_[12]  (.D(\sr_44_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[12]_net_1 ));
    DFN1E1C0 \sr_39_[2]  (.D(\sr_38_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[2]_net_1 ));
    DFN1E1C0 \sr_8_[12]  (.D(\sr_7_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[12]_net_1 ));
    DFN1E1C0 \sr_15_[11]  (.D(\sr_14_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[11]_net_1 ));
    DFN1E1C0 \sr_39_[7]  (.D(\sr_38_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[7]_net_1 ));
    DFN1E1C0 \sr_52_[4]  (.D(\sr_51_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[4]_net_1 ));
    DFN1E1C0 \sr_41_[4]  (.D(\sr_40_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[4]_net_1 ));
    DFN1E1C0 \sr_58_[5]  (.D(\sr_57_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[5]_net_1 ));
    DFN1E1C0 \sr_40_[0]  (.D(\sr_39_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[0]_net_1 ));
    DFN1E1C0 \sr_31_[3]  (.D(\sr_30_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[3]_net_1 ));
    DFN1E1C0 \sr_51_[6]  (.D(\sr_50_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[6]_net_1 ));
    DFN1E1C0 \sr_17_[12]  (.D(\sr_16_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[12]_net_1 ));
    DFN1E1C0 \sr_45_[3]  (.D(\sr_44_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[3]_net_1 ));
    DFN1E1C0 \sr_62_[4]  (.D(\sr_61_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[4]_net_1 ));
    DFN1E1C0 \sr_21_[4]  (.D(\sr_20_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[4]_net_1 ));
    DFN1E1C0 \sr_60_[3]  (.D(\sr_59_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[3]_net_1 ));
    DFN1E1C0 \sr_22_[7]  (.D(\sr_21_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[7]_net_1 ));
    DFN1E1C0 \sr_61_[6]  (.D(\sr_60_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[6]_net_1 ));
    DFN1E1C0 \sr_49_[9]  (.D(\sr_48_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[9]_net_1 ));
    DFN1E1C0 \sr_18_[10]  (.D(\sr_17_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[10]_net_1 ));
    DFN1E1C0 \sr_8_[5]  (.D(\sr_7_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[5]_net_1 ));
    DFN1E1C0 \sr_33_[12]  (.D(\sr_32_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[12]_net_1 ));
    DFN1E1C0 \sr_28_[3]  (.D(\sr_27_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[3]_net_1 ));
    DFN1E1C0 \sr_38_[9]  (.D(\sr_37_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[9]_net_1 ));
    DFN1E1C0 \sr_53_[11]  (.D(\sr_52_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[11]_net_1 ));
    DFN1E1C0 \sr_37_[1]  (.D(\sr_36_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[1]_net_1 ));
    DFN1E1C0 \sr_37_[2]  (.D(\sr_36_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[2]_net_1 ));
    DFN1E1C0 \sr_23_[11]  (.D(\sr_22_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[11]_net_1 ));
    DFN1E1C0 \sr_3_[11]  (.D(\sr_2_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[11]_net_1 ));
    DFN1E1C0 \sr_37_[7]  (.D(\sr_36_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[7]_net_1 ));
    DFN1E1C0 \sr_38_[6]  (.D(\sr_37_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[6]_net_1 ));
    DFN1E1C0 \sr_41_[6]  (.D(\sr_40_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[6]_net_1 ));
    DFN1E1C0 \sr_44_[7]  (.D(\sr_43_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[7]_net_1 ));
    DFN1E1C0 \sr_54_[7]  (.D(\sr_53_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[7]_net_1 ));
    DFN1E1C0 \sr_0_[7]  (.D(cur_error[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[7]));
    DFN1E1C0 \sr_9_[11]  (.D(\sr_8_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[11]_net_1 ));
    DFN1E1C0 \sr_62_[9]  (.D(\sr_61_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[9]_net_1 ));
    DFN1E1C0 \sr_54_[8]  (.D(\sr_53_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[8]_net_1 ));
    DFN1E1C0 \sr_39_[0]  (.D(\sr_38_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[0]_net_1 ));
    DFN1E1C0 \sr_47_[9]  (.D(\sr_46_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[9]_net_1 ));
    DFN1E1C0 \sr_6_[12]  (.D(\sr_5_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[12]_net_1 ));
    DFN1E1C0 \sr_7_[11]  (.D(\sr_6_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[11]_net_1 ));
    DFN1E1C0 \sr_46_[7]  (.D(\sr_45_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[7]_net_1 ));
    DFN1E1C0 \sr_14_[5]  (.D(\sr_13_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[5]_net_1 ));
    DFN1E1C0 \sr_56_[7]  (.D(\sr_55_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[7]_net_1 ));
    DFN1E1C0 \sr_12_[9]  (.D(\sr_11_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[9]_net_1 ));
    DFN1E1C0 \sr_12_[11]  (.D(\sr_11_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[11]_net_1 ));
    DFN1E1C0 \sr_55_[9]  (.D(\sr_54_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[9]_net_1 ));
    DFN1E1C0 \sr_56_[8]  (.D(\sr_55_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[8]_net_1 ));
    DFN1E1C0 \sr_25_[6]  (.D(\sr_24_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[6]_net_1 ));
    DFN1E1C0 \sr_14_[3]  (.D(\sr_13_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[3]_net_1 ));
    DFN1E1C0 \sr_42_[0]  (.D(\sr_41_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[0]_net_1 ));
    DFN1E1C0 \sr_1_[7]  (.D(sr_new[7]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[7]));
    DFN1E1C0 \sr_2_[5]  (.D(sr_prev[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[5]_net_1 ));
    DFN1E1C0 \sr_14_[11]  (.D(\sr_13_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[11]_net_1 ));
    DFN1E1C0 \sr_37_[0]  (.D(\sr_36_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[0]_net_1 ));
    DFN1E1C0 \sr_58_[1]  (.D(\sr_57_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[1]_net_1 ));
    DFN1E1C0 \sr_11_[1]  (.D(\sr_10_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[1]_net_1 ));
    DFN1E1C0 \sr_62_[3]  (.D(\sr_61_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[3]_net_1 ));
    DFN1E1C0 \sr_45_[10]  (.D(\sr_44_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[10]_net_1 ));
    DFN1E1C0 \sr_16_[5]  (.D(\sr_15_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[5]_net_1 ));
    DFN1E1C0 \sr_43_[3]  (.D(\sr_42_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[3]_net_1 ));
    DFN1E1C0 \sr_61_[5]  (.D(\sr_60_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[5]_net_1 ));
    DFN1E1C0 \sr_54_[0]  (.D(\sr_53_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[0]_net_1 ));
    DFN1E1C0 \sr_16_[3]  (.D(\sr_15_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[3]_net_1 ));
    DFN1E1C0 \sr_4_[9]  (.D(\sr_3_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[9]_net_1 ));
    DFN1E1C0 \sr_40_[7]  (.D(\sr_39_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[7]_net_1 ));
    DFN1E1C0 \sr_50_[7]  (.D(\sr_49_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[7]_net_1 ));
    DFN1E1C0 \sr_31_[5]  (.D(\sr_30_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[5]_net_1 ));
    DFN1E1C0 \sr_50_[8]  (.D(\sr_49_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[8]_net_1 ));
    DFN1E1C0 \sr_49_[4]  (.D(\sr_48_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[4]_net_1 ));
    DFN1E1C0 \sr_31_[4]  (.D(\sr_30_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[4]_net_1 ));
    DFN1E1C0 \sr_0_[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable), .Q(sr_new[12]));
    DFN1E1C0 \sr_39_[3]  (.D(\sr_38_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[3]_net_1 ));
    DFN1E1C0 \sr_6_[7]  (.D(\sr_5_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[7]_net_1 ));
    DFN1E1C0 \sr_60_[7]  (.D(\sr_59_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[7]_net_1 ));
    DFN1E1C0 \sr_59_[6]  (.D(\sr_58_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[6]_net_1 ));
    DFN1E1C0 \sr_7_[3]  (.D(\sr_6_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[3]_net_1 ));
    DFN1E1C0 \sr_46_[10]  (.D(\sr_45_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[10]_net_1 ));
    DFN1E1C0 \sr_60_[8]  (.D(\sr_59_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[8]_net_1 ));
    DFN1E1C0 \sr_29_[4]  (.D(\sr_28_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[4]_net_1 ));
    DFN1E1C0 \sr_57_[11]  (.D(\sr_56_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[11]_net_1 ));
    DFN1E1C0 \sr_56_[0]  (.D(\sr_55_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[0]_net_1 ));
    DFN1E1C0 \sr_5_[7]  (.D(\sr_4_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[7]_net_1 ));
    DFN1E1C0 \sr_18_[7]  (.D(\sr_17_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[7]_net_1 ));
    DFN1E1C0 \sr_10_[5]  (.D(\sr_9_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[5]_net_1 ));
    DFN1E1C0 \sr_41_[12]  (.D(\sr_40_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[12]_net_1 ));
    DFN1E1C0 \sr_52_[10]  (.D(\sr_51_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[10]_net_1 ));
    DFN1E1C0 \sr_27_[11]  (.D(\sr_26_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[11]_net_1 ));
    DFN1E1C0 \sr_39_[12]  (.D(\sr_38_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[12]_net_1 ));
    DFN1E1C0 \sr_18_[6]  (.D(\sr_17_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[6]_net_1 ));
    DFN1E1C0 \sr_22_[10]  (.D(\sr_21_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[10]_net_1 ));
    DFN1E1C0 \sr_10_[3]  (.D(\sr_9_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[3]_net_1 ));
    DFN1E1C0 \sr_48_[5]  (.D(\sr_47_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[5]_net_1 ));
    DFN1E1C0 \sr_60_[0]  (.D(\sr_59_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[0]_net_1 ));
    DFN1E1C0 \sr_47_[4]  (.D(\sr_46_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[4]_net_1 ));
    DFN1E1C0 \sr_30_[12]  (.D(\sr_29_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[12]_net_1 ));
    DFN1E1C0 \sr_37_[3]  (.D(\sr_36_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[3]_net_1 ));
    DFN1E1C0 \sr_57_[6]  (.D(\sr_56_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[6]_net_1 ));
    DFN1E1C0 \sr_49_[6]  (.D(\sr_48_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[6]_net_1 ));
    DFN1E1C0 \sr_3_[3]  (.D(\sr_2_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[3]_net_1 ));
    DFN1E1C0 \sr_28_[9]  (.D(\sr_27_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[9]_net_1 ));
    DFN1E1C0 \sr_27_[4]  (.D(\sr_26_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[4]_net_1 ));
    DFN1E1C0 \sr_62_[12]  (.D(\sr_61_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[12]_net_1 ));
    DFN1E1C0 \sr_50_[0]  (.D(\sr_49_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[0]_net_1 ));
    DFN1E1C0 \sr_53_[9]  (.D(\sr_52_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[9]_net_1 ));
    DFN1E1C0 \sr_23_[6]  (.D(\sr_22_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[6]_net_1 ));
    DFN1E1C0 \sr_28_[1]  (.D(\sr_27_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[1]_net_1 ));
    DFN1E1C0 \sr_11_[4]  (.D(\sr_10_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[4]_net_1 ));
    DFN1E1C0 \sr_30_[10]  (.D(\sr_29_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[10]_net_1 ));
    DFN1E1C0 \sr_21_[8]  (.D(\sr_20_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[8]_net_1 ));
    DFN1E1C0 \sr_16_[12]  (.D(\sr_15_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[12]_net_1 ));
    DFN1E1C0 \sr_41_[10]  (.D(\sr_40_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[10]_net_1 ));
    DFN1E1C0 \sr_45_[1]  (.D(\sr_44_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[1]_net_1 ));
    DFN1E1C0 \sr_33_[10]  (.D(\sr_32_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[10]_net_1 ));
    DFN1E1C0 \sr_14_[12]  (.D(\sr_13_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[12]_net_1 ));
    DFN1E1C0 \sr_41_[11]  (.D(\sr_40_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[11]_net_1 ));
    DFN1E1C0 \sr_55_[12]  (.D(\sr_54_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[12]_net_1 ));
    DFN1E1C0 \sr_42_[7]  (.D(\sr_41_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[7]_net_1 ));
    DFN1E1C0 \sr_52_[7]  (.D(\sr_51_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[7]_net_1 ));
    DFN1E1C0 \sr_41_[2]  (.D(\sr_40_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[2]_net_1 ));
    DFN1E1C0 \sr_52_[8]  (.D(\sr_51_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[8]_net_1 ));
    DFN1E1C0 \sr_25_[12]  (.D(\sr_24_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[12]_net_1 ));
    DFN1E1C0 \sr_47_[6]  (.D(\sr_46_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[6]_net_1 ));
    DFN1E1C0 \sr_62_[7]  (.D(\sr_61_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[7]_net_1 ));
    DFN1E1C0 \sr_62_[8]  (.D(\sr_61_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[8]_net_1 ));
    DFN1E1C0 \sr_19_[1]  (.D(\sr_18_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[1]_net_1 ));
    DFN1E1C0 \sr_21_[0]  (.D(\sr_20_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[0]_net_1 ));
    DFN1E1C0 \sr_39_[10]  (.D(\sr_38_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[10]_net_1 ));
    DFN1E1C0 \sr_12_[5]  (.D(\sr_11_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[5]_net_1 ));
    DFN1E1C0 \sr_0_[10]  (.D(cur_error[10]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable), .Q(sr_new[10]));
    DFN1E1C0 \sr_12_[3]  (.D(\sr_11_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[3]_net_1 ));
    DFN1E1C0 \sr_34_[1]  (.D(\sr_33_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[1]_net_1 ));
    DFN1E1C0 \sr_39_[5]  (.D(\sr_38_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[5]_net_1 ));
    DFN1E1C0 \sr_5_[11]  (.D(\sr_4_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[11]_net_1 ));
    DFN1E1C0 \sr_34_[2]  (.D(\sr_33_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[2]_net_1 ));
    DFN1E1C0 \sr_39_[4]  (.D(\sr_38_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[4]_net_1 ));
    DFN1E1C0 \sr_55_[2]  (.D(\sr_54_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[2]_net_1 ));
    DFN1E1C0 \sr_62_[0]  (.D(\sr_61_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[0]_net_1 ));
    DFN1E1C0 \sr_34_[7]  (.D(\sr_33_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[7]_net_1 ));
    DFN1E1C0 \sr_41_[8]  (.D(\sr_40_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[8]_net_1 ));
    DFN1E1C0 \sr_52_[0]  (.D(\sr_51_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[0]_net_1 ));
    DFN1E1C0 \sr_17_[1]  (.D(\sr_16_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[1]_net_1 ));
    DFN1E1C0 \sr_4_[0]  (.D(\sr_3_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[0]_net_1 ));
    DFN1E1C0 \sr_36_[1]  (.D(\sr_35_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[1]_net_1 ));
    DFN1E1C0 \sr_13_[12]  (.D(\sr_12_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[12]_net_1 ));
    DFN1E1C0 \sr_4_[6]  (.D(\sr_3_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[6]_net_1 ));
    DFN1E1C0 \sr_44_[9]  (.D(\sr_43_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[9]_net_1 ));
    DFN1E1C0 \sr_0_[3]  (.D(cur_error[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[3]));
    DFN1E1C0 \sr_36_[2]  (.D(\sr_35_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[2]_net_1 ));
    DFN1E1C0 \sr_51_[3]  (.D(\sr_50_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[3]_net_1 ));
    DFN1E1C0 \sr_36_[7]  (.D(\sr_35_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[7]_net_1 ));
    DFN1E1C0 \sr_21_[2]  (.D(\sr_20_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[2]_net_1 ));
    DFN1E1C0 \sr_37_[5]  (.D(\sr_36_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[5]_net_1 ));
    DFN1E1C0 \sr_55_[4]  (.D(\sr_54_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[4]_net_1 ));
    DFN1E1C0 \sr_21_[5]  (.D(\sr_20_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[5]_net_1 ));
    DFN1E1C0 \sr_43_[1]  (.D(\sr_42_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[1]_net_1 ));
    DFN1E1C0 \sr_11_[8]  (.D(\sr_10_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[8]_net_1 ));
    DFN1E1C0 \sr_37_[4]  (.D(\sr_36_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[4]_net_1 ));
    DFN1E1C0 \sr_62_[11]  (.D(\sr_61_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[11]_net_1 ));
    DFN1E1C0 \sr_46_[9]  (.D(\sr_45_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[9]_net_1 ));
    DFN1E1C0 \sr_25_[7]  (.D(\sr_24_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[7]_net_1 ));
    DFN1E1C0 \sr_48_[3]  (.D(\sr_47_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[3]_net_1 ));
    DFN1E1C0 \sr_30_[1]  (.D(\sr_29_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[1]_net_1 ));
    DFN1E1C0 \sr_4_[1]  (.D(\sr_3_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[1]_net_1 ));
    DFN1E1C0 \sr_55_[10]  (.D(\sr_54_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[10]_net_1 ));
    DFN1E1C0 \sr_19_[4]  (.D(\sr_18_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[4]_net_1 ));
    DFN1E1C0 \sr_9_[7]  (.D(\sr_8_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[7]_net_1 ));
    DFN1E1C0 \sr_7_[4]  (.D(\sr_6_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[4]_net_1 ));
    DFN1E1C0 \sr_29_[8]  (.D(\sr_28_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[8]_net_1 ));
    DFN1E1C0 \sr_1_[3]  (.D(sr_new[3]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[3]));
    DFN1E1C0 \sr_34_[0]  (.D(\sr_33_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[0]_net_1 ));
    DFN1E1C0 \sr_30_[2]  (.D(\sr_29_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[2]_net_1 ));
    DFN1E1C0 \sr_25_[10]  (.D(\sr_24_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[10]_net_1 ));
    DFN1E1C0 \sr_30_[7]  (.D(\sr_29_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[7]_net_1 ));
    DFN1E1C0 \sr_49_[2]  (.D(\sr_48_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[2]_net_1 ));
    DFN1E1C0 \sr_56_[10]  (.D(\sr_55_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[10]_net_1 ));
    DFN1E1C0 \sr_40_[9]  (.D(\sr_39_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[9]_net_1 ));
    DFN1E1C0 \sr_36_[0]  (.D(\sr_35_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[0]_net_1 ));
    DFN1E1C0 \sr_11_[2]  (.D(\sr_10_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[2]_net_1 ));
    DFN1E1C0 \sr_30_[11]  (.D(\sr_29_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[11]_net_1 ));
    DFN1E1C0 \sr_53_[2]  (.D(\sr_52_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[2]_net_1 ));
    DFN1E1C0 \sr_26_[10]  (.D(\sr_25_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[10]_net_1 ));
    DFN1E1C0 \sr_11_[0]  (.D(\sr_10_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[0]_net_1 ));
    DFN1E1C0 \sr_31_[8]  (.D(\sr_30_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[8]_net_1 ));
    DFN1E1C0 \sr_29_[0]  (.D(\sr_28_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[0]_net_1 ));
    DFN1E1C0 \sr_17_[4]  (.D(\sr_16_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[4]_net_1 ));
    DFN1E1C0 \sr_6_[3]  (.D(\sr_5_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[3]_net_1 ));
    DFN1E1C0 \sr_51_[12]  (.D(\sr_50_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[12]_net_1 ));
    DFN1E1C0 \sr_27_[8]  (.D(\sr_26_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[8]_net_1 ));
    DFN1E1C0 \sr_3_[4]  (.D(\sr_2_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[4]_net_1 ));
    DFN1E1C0 \sr_63_[2]  (.D(\sr_62_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[2]));
    DFN1E1C0 \sr_21_[12]  (.D(\sr_20_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[12]_net_1 ));
    DFN1E1C0 \sr_5_[3]  (.D(\sr_4_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[3]_net_1 ));
    DFN1E1C0 \sr_15_[9]  (.D(\sr_14_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[9]_net_1 ));
    DFN1E1C0 \sr_51_[5]  (.D(\sr_50_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[5]_net_1 ));
    DFN1E1C0 \sr_47_[2]  (.D(\sr_46_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[2]_net_1 ));
    DFN1E1C0 \sr_47_[10]  (.D(\sr_46_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[10]_net_1 ));
    DFN1E1C0 \sr_45_[0]  (.D(\sr_44_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[0]_net_1 ));
    DFN1E1C0 \sr_58_[9]  (.D(\sr_57_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[9]_net_1 ));
    DFN1E1C0 \sr_30_[0]  (.D(\sr_29_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[0]_net_1 ));
    DFN1E1C0 \sr_44_[4]  (.D(\sr_43_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[4]_net_1 ));
    DFN1E1C0 \sr_53_[4]  (.D(\sr_52_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[4]_net_1 ));
    DFN1E1C0 \sr_34_[3]  (.D(\sr_33_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[3]_net_1 ));
    DFN1E1C0 \sr_54_[6]  (.D(\sr_53_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[6]_net_1 ));
    DFN1E1C0 \sr_49_[8]  (.D(\sr_48_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[8]_net_1 ));
    DFN1E1C0 \sr_28_[6]  (.D(\sr_27_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[6]_net_1 ));
    DFN1E1C0 \sr_21_[3]  (.D(\sr_20_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[3]_net_1 ));
    DFN1E1C0 \sr_31_[9]  (.D(\sr_30_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[9]_net_1 ));
    DFN1E1C0 \sr_8_[7]  (.D(\sr_7_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[7]_net_1 ));
    DFN1E1C0 \sr_27_[0]  (.D(\sr_26_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[0]_net_1 ));
    DFN1E1C0 \sr_24_[4]  (.D(\sr_23_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[4]_net_1 ));
    DFN1E1C0 \sr_63_[4]  (.D(\sr_62_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[4]));
    DFN1E1C0 \sr_32_[1]  (.D(\sr_31_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[1]_net_1 ));
    DFN1E1C0 \sr_19_[12]  (.D(\sr_18_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[12]_net_1 ));
    DFN1E1C0 \sr_23_[7]  (.D(\sr_22_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[7]_net_1 ));
    DFN1E1C0 \sr_51_[10]  (.D(\sr_50_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[10]_net_1 ));
    DFN1E1C0 \sr_32_[2]  (.D(\sr_31_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[2]_net_1 ));
    DFN1E1C0 \sr_38_[12]  (.D(\sr_37_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[12]_net_1 ));
    DFN1E1C0 \sr_59_[3]  (.D(\sr_58_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[3]_net_1 ));
    DFN1E1C0 \sr_51_[11]  (.D(\sr_50_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[11]_net_1 ));
    DFN1E1C0 \sr_29_[2]  (.D(\sr_28_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[2]_net_1 ));
    DFN1E1C0 \sr_32_[7]  (.D(\sr_31_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[7]_net_1 ));
    DFN1E1C0 \sr_21_[10]  (.D(\sr_20_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[10]_net_1 ));
    DFN1E1C0 \sr_46_[4]  (.D(\sr_45_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[4]_net_1 ));
    DFN1E1C0 \sr_31_[6]  (.D(\sr_30_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[6]_net_1 ));
    DFN1E1C0 \sr_36_[3]  (.D(\sr_35_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[3]_net_1 ));
    DFN1E1C0 \sr_29_[5]  (.D(\sr_28_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[5]_net_1 ));
    DFN1E1C0 \sr_56_[6]  (.D(\sr_55_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[6]_net_1 ));
    DFN1E1C0 \sr_21_[11]  (.D(\sr_20_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[11]_net_1 ));
    DFN1E1C0 \sr_19_[8]  (.D(\sr_18_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[8]_net_1 ));
    DFN1E1C0 \sr_44_[10]  (.D(\sr_43_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[10]_net_1 ));
    DFN1E1C0 \sr_10_[12]  (.D(\sr_9_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[12]_net_1 ));
    DFN1E1C0 \sr_26_[4]  (.D(\sr_25_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[4]_net_1 ));
    DFN1E1C0 \sr_47_[8]  (.D(\sr_46_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[8]_net_1 ));
    DFN1E1C0 \sr_44_[6]  (.D(\sr_43_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[6]_net_1 ));
    DFN1E1C0 \sr_42_[9]  (.D(\sr_41_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[9]_net_1 ));
    DFN1E1C0 \sr_63_[9]  (.D(\sr_62_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[9]));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \sr_10_[10]  (.D(\sr_9_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[10]_net_1 ));
    DFN1E1C0 \sr_2_[10]  (.D(sr_prev[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[10]_net_1 ));
    DFN1E1C0 \sr_13_[10]  (.D(\sr_12_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[10]_net_1 ));
    DFN1E1C0 \sr_57_[3]  (.D(\sr_56_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[3]_net_1 ));
    DFN1E1C0 \sr_27_[2]  (.D(\sr_26_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[2]_net_1 ));
    DFN1E1C0 \sr_40_[4]  (.D(\sr_39_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[4]_net_1 ));
    DFN1E1C0 \sr_30_[3]  (.D(\sr_29_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[3]_net_1 ));
    DFN1E1C0 \sr_50_[6]  (.D(\sr_49_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[6]_net_1 ));
    DFN1E1C0 \sr_27_[5]  (.D(\sr_26_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[5]_net_1 ));
    DFN1E1C0 \sr_46_[6]  (.D(\sr_45_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[6]_net_1 ));
    DFN1E1C0 \sr_38_[11]  (.D(\sr_37_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[11]_net_1 ));
    DFN1E1C0 \sr_17_[8]  (.D(\sr_16_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[8]_net_1 ));
    DFN1E1C0 \sr_20_[4]  (.D(\sr_19_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[4]_net_1 ));
    DFN1E1C0 \sr_0_[4]  (.D(cur_error[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[4]));
    DFN1E1C0 \sr_49_[11]  (.D(\sr_48_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[11]_net_1 ));
    DFN1E1C0 \sr_13_[9]  (.D(\sr_12_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[9]_net_1 ));
    DFN1E1C0 \sr_60_[6]  (.D(\sr_59_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[6]_net_1 ));
    DFN1E1C0 \sr_2_[7]  (.D(sr_prev[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[7]_net_1 ));
    DFN1E1C0 \sr_51_[1]  (.D(\sr_50_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[1]_net_1 ));
    DFN1E1C0 \sr_32_[0]  (.D(\sr_31_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[0]_net_1 ));
    DFN1E1C0 \sr_7_[2]  (.D(\sr_6_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[2]_net_1 ));
    DFN1E1C0 \sr_4_[11]  (.D(\sr_3_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[11]_net_1 ));
    DFN1E1C0 \sr_19_[2]  (.D(\sr_18_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[2]_net_1 ));
    DFN1E1C0 \sr_7_[8]  (.D(\sr_6_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[8]_net_1 ));
    DFN1E1C0 \sr_4_[5]  (.D(\sr_3_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[5]_net_1 ));
    DFN1E1C0 \sr_43_[0]  (.D(\sr_42_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[0]_net_1 ));
    DFN1E1C0 \sr_19_[0]  (.D(\sr_18_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[0]_net_1 ));
    DFN1E1C0 \sr_9_[10]  (.D(\sr_8_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[10]_net_1 ));
    DFN1E1C0 \sr_39_[8]  (.D(\sr_38_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[8]_net_1 ));
    DFN1E1C0 \sr_61_[1]  (.D(\sr_60_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[1]_net_1 ));
    DFN1E1C0 \sr_19_[10]  (.D(\sr_18_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[10]_net_1 ));
    DFN1E1C0 \sr_14_[1]  (.D(\sr_13_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[1]_net_1 ));
    DFN1E1C0 \sr_63_[3]  (.D(\sr_62_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[3]));
    DFN1E1C0 \sr_45_[7]  (.D(\sr_44_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[7]_net_1 ));
    DFN1E1C0 \sr_59_[5]  (.D(\sr_58_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[5]_net_1 ));
    DFN1E1C0 \sr_55_[7]  (.D(\sr_54_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[7]_net_1 ));
    DFN1E1C0 \sr_63_[12]  (.D(\sr_62_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[12]));
    DFN1E1C0 \sr_48_[1]  (.D(\sr_47_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[1]_net_1 ));
    DFN1E1C0 \sr_42_[12]  (.D(\sr_41_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[12]_net_1 ));
    DFN1E1C0 \sr_40_[6]  (.D(\sr_39_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[6]_net_1 ));
    DFN1E1C0 \sr_55_[8]  (.D(\sr_54_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[8]_net_1 ));
    DFN1E1C0 \sr_1_[4]  (.D(sr_new[4]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[4]));
    DFN1E1C0 \sr_34_[5]  (.D(\sr_33_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[5]_net_1 ));
    DFN1E1C0 \sr_6_[11]  (.D(\sr_5_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[11]_net_1 ));
    DFN1E1C0 \sr_11_[7]  (.D(\sr_10_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[7]_net_1 ));
    DFN1E1C0 \sr_34_[4]  (.D(\sr_33_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[4]_net_1 ));
    DFN1E1C0 \sr_16_[1]  (.D(\sr_15_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[1]_net_1 ));
    DFN1E1C0 \sr_29_[3]  (.D(\sr_28_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[3]_net_1 ));
    DFN1E1C0 \sr_17_[2]  (.D(\sr_16_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[2]_net_1 ));
    DFN1E1C0 \sr_39_[9]  (.D(\sr_38_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[9]_net_1 ));
    DFN1E1C0 \sr_3_[2]  (.D(\sr_2_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[2]_net_1 ));
    DFN1E1C0 \sr_46_[11]  (.D(\sr_45_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[11]_net_1 ));
    DFN1E1C0 \sr_3_[8]  (.D(\sr_2_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[8]_net_1 ));
    DFN1E1C0 \sr_33_[11]  (.D(\sr_32_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[11]_net_1 ));
    DFN1E1C0 \sr_17_[0]  (.D(\sr_16_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[0]_net_1 ));
    DFN1E1C0 \sr_37_[8]  (.D(\sr_36_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[8]_net_1 ));
    DFN1E1C0 \sr_15_[5]  (.D(\sr_14_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[5]_net_1 ));
    DFN1E1C0 \sr_11_[6]  (.D(\sr_10_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[6]_net_1 ));
    
endmodule


module controller_Z1_4(
       state_0_d0,
       state_0_0,
       pwm_chg,
       sig_prev_0,
       sig_old_i_0_0,
       N_46_1,
       avg_done,
       sig_old_i_0,
       sig_prev,
       sum_rdy,
       deriv_enable,
       calc_avg,
       calc_int,
       pwm_enable,
       sum_enable,
       calc_error,
       avg_enable,
       int_enable,
       pwm_chg_0,
       avg_enable_0,
       n_rst_c,
       clk_c,
       avg_enable_1
    );
input  state_0_d0;
input  state_0_0;
output pwm_chg;
input  sig_prev_0;
input  sig_old_i_0_0;
input  N_46_1;
input  avg_done;
input  sig_old_i_0;
input  sig_prev;
input  sum_rdy;
output deriv_enable;
output calc_avg;
output calc_int;
output pwm_enable;
output sum_enable;
output calc_error;
output avg_enable;
output int_enable;
output pwm_chg_0;
output avg_enable_0;
input  n_rst_c;
input  clk_c;
output avg_enable_1;

    wire \state_RNIKCLT1[0]_net_1 , N_12, \state[5]_net_1 , N_94, 
        count_31_0, count_c13, count_n14, \count[14]_net_1 , N_62, 
        count_n13, count_c12, \count[13]_net_1 , count_n12, count_c11, 
        \count[12]_net_1 , count_n15, \count[15]_net_1 , count_c7, 
        count_c6, \count[7]_net_1 , count_c5, \count[6]_net_1 , 
        count_c4, \count[5]_net_1 , count_c3, \count[4]_net_1 , 
        count_c2, \count[3]_net_1 , \count[1]_net_1 , \count[0]_net_1 , 
        \count[2]_net_1 , count_c8, \count[8]_net_1 , count_c9, 
        \count[9]_net_1 , count_c10, \count[10]_net_1 , 
        \count[11]_net_1 , \state_ns_0_a2_9[0] , \state[10]_net_1 , 
        N_33, \state_ns_0_a2_8[0] , \state_ns_0_a2_6[0] , 
        \state_ns_0_a2_5[0] , \state_ns_0_a2_2[0] , N_270, N_272, 
        \state_ns_0_a2_1[0] , \state_ns_0_a2_0[0] , \state[7]_net_1 , 
        next_state_0_sqmuxa_1_1_a2_0_a2_0, \state_ns_i_0_0[2] , 
        un1_countlto15_13, un1_countlto15_5, un1_countlto15_4, 
        un1_countlto15_11, un1_countlto15_12, un1_countlto15_1, 
        un1_countlto15_0, un1_countlto15_9, un1_countlto15_7, 
        un1_countlto15_3, N_274, N_23, N_273, \state[0]_net_1 , N_26, 
        next_state15_li, \state_RNIL4T11[4]_net_1 , 
        \state_RNO[5]_net_1 , N_24, count_n7, count_n6, count_n5, 
        count_n4, count_n3, count_n2, count_n2_tz, count_n8, count_n9, 
        count_n10, count_n11, \state_ns[4] , \state[4]_net_1 , 
        \state_RNO[8]_net_1 , \state[12]_net_1 , \state_ns[10] , 
        \state_ns[0] , \state_ns[1] , \avg_count[1]_net_1 , 
        \avg_count[0]_net_1 , \state_ns[7] , \state_ns[12] , N_27, 
        count_n1, N_267, counte, \DWACT_ADD_CI_0_partial_sum[0] , I_10, 
        \DWACT_ADD_CI_0_TMP[0] , GND, VCC;
    
    OR2B \state_RNI7D0A[12]  (.A(\state[12]_net_1 ), .B(
        \state[4]_net_1 ), .Y(N_273));
    NOR3C \count_RNINV863[7]  (.A(un1_countlto15_5), .B(
        un1_countlto15_4), .C(un1_countlto15_11), .Y(un1_countlto15_13)
        );
    DFN1E1C0 \count[5]  (.D(count_n5), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[5]_net_1 ));
    OA1A \state_RNO_0[0]  (.A(\state[10]_net_1 ), .B(N_33), .C(
        \state_ns_0_a2_8[0] ), .Y(\state_ns_0_a2_9[0] ));
    DFN1E1C0 \count[1]  (.D(count_n1), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[1]_net_1 ));
    NOR2B \count_RNISOSK2[7]  (.A(count_c6), .B(\count[7]_net_1 ), .Y(
        count_c7));
    NOR2B \count_RNI529A2[6]  (.A(count_c5), .B(\count[6]_net_1 ), .Y(
        count_c6));
    DFN1E1C0 \count[10]  (.D(count_n10), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[10]_net_1 ));
    DFN1E1C0 \count[0]  (.D(N_267), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[0]_net_1 ));
    NOR2 \state_RNO_9[0]  (.A(calc_avg), .B(deriv_enable), .Y(
        \state_ns_0_a2_0[0] ));
    DFN1C0 \state[13]  (.D(N_12), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_chg));
    DFN1E1C0 \count[14]  (.D(count_n14), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[14]_net_1 ));
    NOR2 \count_RNIBA7L[5]  (.A(\count[6]_net_1 ), .B(\count[5]_net_1 )
        , .Y(un1_countlto15_3));
    DFN1C0 \state[7]  (.D(\state_ns[7] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[7]_net_1 ));
    NOR2 \state_RNIFHUF[0]  (.A(\state[0]_net_1 ), .B(N_272), .Y(N_23));
    DFN1C0 \state[5]  (.D(\state_RNO[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[5]_net_1 ));
    XA1B \count_RNO[7]  (.A(\count[7]_net_1 ), .B(count_c6), .C(N_62), 
        .Y(count_n7));
    AX1 \count_RNO[15]  (.A(N_62), .B(\count[15]_net_1 ), .C(N_94), .Y(
        count_n15));
    NOR3C \count_RNIBTBO2[2]  (.A(un1_countlto15_1), .B(
        un1_countlto15_0), .C(un1_countlto15_9), .Y(un1_countlto15_12));
    AO1 \state_RNIEAMV6[10]  (.A(sig_old_i_0_0), .B(sig_prev_0), .C(
        N_62), .Y(counte));
    DFN1C0 \state[4]  (.D(\state_ns[4] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[4]_net_1 ));
    NOR2A \count_RNO[2]  (.A(count_n2_tz), .B(N_62), .Y(count_n2));
    AO1A \state_RNO[7]  (.A(N_46_1), .B(\state[7]_net_1 ), .C(calc_int)
        , .Y(\state_ns[7] ));
    DFN1C0 \state_1[2]  (.D(\state_RNIKCLT1[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable_1));
    NOR2B \count_RNIJECK4[12]  (.A(count_c11), .B(\count[12]_net_1 ), 
        .Y(count_c12));
    NOR2A \state_RNO_0[5]  (.A(N_272), .B(\state[10]_net_1 ), .Y(N_24));
    DFN1C0 \state_0[2]  (.D(\state_RNIKCLT1[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable_0));
    XA1B \count_RNO[9]  (.A(count_c8), .B(\count[9]_net_1 ), .C(N_62), 
        .Y(count_n9));
    DFN1C0 \state[6]  (.D(int_enable), .CLK(clk_c), .CLR(n_rst_c), .Q(
        calc_int));
    NOR2 \state_RNO_6[0]  (.A(sum_enable), .B(\state[7]_net_1 ), .Y(
        \state_ns_0_a2_2[0] ));
    DFN1C0 \state[2]  (.D(\state_RNIKCLT1[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable));
    NOR3A \count_RNIE2BO1[11]  (.A(un1_countlto15_7), .B(
        \count[12]_net_1 ), .C(\count[11]_net_1 ), .Y(
        un1_countlto15_11));
    VCC VCC_i (.Y(VCC));
    XOR2 un1_avg_count_1_I_10 (.A(\avg_count[1]_net_1 ), .B(
        \DWACT_ADD_CI_0_TMP[0] ), .Y(I_10));
    NOR2B \count_RNIKGGV2[8]  (.A(count_c7), .B(\count[8]_net_1 ), .Y(
        count_c8));
    NOR3A \count_RNIIGEA1[3]  (.A(un1_countlto15_3), .B(
        \count[3]_net_1 ), .C(\count[4]_net_1 ), .Y(un1_countlto15_9));
    XA1B \count_RNO[4]  (.A(\count[4]_net_1 ), .B(count_c3), .C(N_62), 
        .Y(count_n4));
    DFN1C0 \state[3]  (.D(avg_enable), .CLK(clk_c), .CLR(n_rst_c), .Q(
        calc_avg));
    NOR2B \count_RNI64EA1[3]  (.A(count_c2), .B(\count[3]_net_1 ), .Y(
        count_c3));
    DFN1E1C0 \count[8]  (.D(count_n8), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[8]_net_1 ));
    OR2B \avg_count_RNIRD3J[1]  (.A(\avg_count[1]_net_1 ), .B(
        \avg_count[0]_net_1 ), .Y(next_state15_li));
    NOR3 \state_RNIKCLT1[0]  (.A(N_274), .B(\state_ns_i_0_0[2] ), .C(
        N_23), .Y(\state_RNIKCLT1[0]_net_1 ));
    NOR2B \state_RNIIBHB[10]  (.A(\state[10]_net_1 ), .B(sum_rdy), .Y(
        next_state_0_sqmuxa_1_1_a2_0_a2_0));
    XA1B \count_RNO[10]  (.A(count_c9), .B(\count[10]_net_1 ), .C(N_62)
        , .Y(count_n10));
    NOR2B \state_RNO[8]  (.A(\state[7]_net_1 ), .B(N_46_1), .Y(
        \state_RNO[8]_net_1 ));
    NOR2B \state_RNIL4T11[4]  (.A(\state[4]_net_1 ), .B(avg_done), .Y(
        \state_RNIL4T11[4]_net_1 ));
    NOR2B \count_RNIQN1L1[4]  (.A(count_c3), .B(\count[4]_net_1 ), .Y(
        count_c4));
    NOR3B \state_RNO_1[0]  (.A(next_state15_li), .B(
        \state_RNIL4T11[4]_net_1 ), .C(\state[10]_net_1 ), .Y(N_26));
    AOI1B \state_RNIK86A6[10]  (.A(un1_countlto15_13), .B(
        un1_countlto15_12), .C(next_state_0_sqmuxa_1_1_a2_0_a2_0), .Y(
        N_62));
    CLKINT \state_RNID9U5[5]  (.A(\state[5]_net_1 ), .Y(int_enable));
    DFN1E1C0 \count[15]  (.D(count_n15), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[15]_net_1 ));
    XA1B \count_RNO[3]  (.A(\count[3]_net_1 ), .B(count_c2), .C(N_62), 
        .Y(count_n3));
    NOR3C \count_RNIJHQV[2]  (.A(\count[1]_net_1 ), .B(
        \count[0]_net_1 ), .C(\count[2]_net_1 ), .Y(count_c2));
    DFN1E1C0 \count[11]  (.D(count_n11), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[11]_net_1 ));
    OA1 \state_RNO_0[12]  (.A(state_0_0), .B(state_0_d0), .C(
        \state[12]_net_1 ), .Y(N_27));
    DFN1C0 \state_0[13]  (.D(N_12), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_chg_0));
    XA1B \count_RNO[8]  (.A(count_c7), .B(\count[8]_net_1 ), .C(N_62), 
        .Y(count_n8));
    OR2 \state_RNI7D0A_0[12]  (.A(\state[12]_net_1 ), .B(
        \state[4]_net_1 ), .Y(N_272));
    AO1A \state_RNO[10]  (.A(sum_rdy), .B(\state[10]_net_1 ), .C(
        sum_enable), .Y(\state_ns[10] ));
    DFN1E1C0 \count[13]  (.D(count_n13), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[13]_net_1 ));
    XA1B \count_RNO[5]  (.A(\count[5]_net_1 ), .B(count_c4), .C(N_62), 
        .Y(count_n5));
    XA1B \count_RNO[1]  (.A(\count[1]_net_1 ), .B(\count[0]_net_1 ), 
        .C(N_62), .Y(count_n1));
    XA1B \count_RNO[11]  (.A(count_c10), .B(\count[11]_net_1 ), .C(
        N_62), .Y(count_n11));
    NOR2B \count_RNIEV6O3[10]  (.A(count_c9), .B(\count[10]_net_1 ), 
        .Y(count_c10));
    NOR3B \state_RNO_4[0]  (.A(\state_ns_0_a2_2[0] ), .B(N_270), .C(
        N_272), .Y(\state_ns_0_a2_6[0] ));
    DFN1C0 \state[11]  (.D(N_62), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_enable));
    DFN1E1C0 \count[2]  (.D(count_n2), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[2]_net_1 ));
    DFN1P0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .PRE(n_rst_c), 
        .Q(\state[0]_net_1 ));
    NOR2B \count_RNIFCLV1[5]  (.A(count_c4), .B(\count[5]_net_1 ), .Y(
        count_c5));
    NOR2 \count_RNIFE7L[7]  (.A(\count[7]_net_1 ), .B(\count[8]_net_1 )
        , .Y(un1_countlto15_4));
    NOR3A \state_RNI8K0K[0]  (.A(N_273), .B(\state[10]_net_1 ), .C(
        \state[0]_net_1 ), .Y(N_274));
    DFN1C0 \state[12]  (.D(\state_ns[12] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[12]_net_1 ));
    NOR2A \count_RNO_1[15]  (.A(\count[14]_net_1 ), .B(N_62), .Y(
        count_31_0));
    NOR2 \count_RNIQEMO[9]  (.A(\count[9]_net_1 ), .B(
        \count[10]_net_1 ), .Y(un1_countlto15_5));
    GND GND_i (.Y(GND));
    NOR2 \count_RNI327L[2]  (.A(\count[2]_net_1 ), .B(\count[1]_net_1 )
        , .Y(un1_countlto15_1));
    DFN1E1C0 \count[9]  (.D(count_n9), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[9]_net_1 ));
    XA1B \count_RNO[6]  (.A(\count[6]_net_1 ), .B(count_c5), .C(N_62), 
        .Y(count_n6));
    XA1B \count_RNO[12]  (.A(count_c11), .B(\count[12]_net_1 ), .C(
        N_62), .Y(count_n12));
    NOR2 \count_RNO[0]  (.A(\count[0]_net_1 ), .B(N_62), .Y(N_267));
    AND2 un1_avg_count_1_I_1 (.A(\avg_count[0]_net_1 ), .B(
        \state_RNIL4T11[4]_net_1 ), .Y(\DWACT_ADD_CI_0_TMP[0] ));
    XOR2 un1_avg_count_1_I_8 (.A(\avg_count[0]_net_1 ), .B(
        \state_RNIL4T11[4]_net_1 ), .Y(\DWACT_ADD_CI_0_partial_sum[0] )
        );
    NOR2B \count_RNIN7F25[13]  (.A(count_c12), .B(\count[13]_net_1 ), 
        .Y(count_c13));
    NOR2 \count_RNI9J5S[13]  (.A(\count[14]_net_1 ), .B(
        \count[13]_net_1 ), .Y(un1_countlto15_7));
    NOR3B \state_RNO_5[0]  (.A(\state_ns_0_a2_1[0] ), .B(
        \state_ns_0_a2_0[0] ), .C(calc_error), .Y(\state_ns_0_a2_5[0] )
        );
    NOR3C \state_RNO_2[0]  (.A(un1_countlto15_12), .B(
        un1_countlto15_13), .C(sum_rdy), .Y(N_33));
    AO1A \state_RNO[4]  (.A(avg_done), .B(\state[4]_net_1 ), .C(
        calc_avg), .Y(\state_ns[4] ));
    DFN1E1C0 \count[6]  (.D(count_n6), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[6]_net_1 ));
    OR2 \state_RNO[12]  (.A(N_27), .B(pwm_enable), .Y(\state_ns[12] ));
    DFN1C0 \state[10]  (.D(\state_ns[10] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[10]_net_1 ));
    DFN1E1C0 \count[3]  (.D(count_n3), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[3]_net_1 ));
    DFN1C0 \state[1]  (.D(\state_ns[1] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(calc_error));
    NOR2 \state_RNO_8[0]  (.A(pwm_enable), .B(calc_int), .Y(
        \state_ns_0_a2_1[0] ));
    DFN1C0 \state[8]  (.D(\state_RNO[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(deriv_enable));
    NOR2B \count_RNIGM964[11]  (.A(count_c10), .B(\count[11]_net_1 ), 
        .Y(count_c11));
    AX1C \count_RNO_0[2]  (.A(\count[1]_net_1 ), .B(\count[0]_net_1 ), 
        .C(\count[2]_net_1 ), .Y(count_n2_tz));
    NOR3A \state_RNO[5]  (.A(calc_error), .B(\state[7]_net_1 ), .C(
        N_24), .Y(\state_RNO[5]_net_1 ));
    XA1B \count_RNO[14]  (.A(count_c13), .B(\count[14]_net_1 ), .C(
        N_62), .Y(count_n14));
    NOR2 \count_RNIMAMO[15]  (.A(\count[15]_net_1 ), .B(
        \count[0]_net_1 ), .Y(un1_countlto15_0));
    XA1B \count_RNO[13]  (.A(count_c12), .B(\count[13]_net_1 ), .C(
        N_62), .Y(count_n13));
    DFN1C0 \state[9]  (.D(deriv_enable), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(sum_enable));
    NOR3A \state_RNIGBH9[12]  (.A(\state[12]_net_1 ), .B(state_0_0), 
        .C(state_0_d0), .Y(N_12));
    NOR2B \count_RNID94A3[9]  (.A(count_c8), .B(\count[9]_net_1 ), .Y(
        count_c9));
    DFN1C0 \avg_count[0]  (.D(\DWACT_ADD_CI_0_partial_sum[0] ), .CLK(
        clk_c), .CLR(n_rst_c), .Q(\avg_count[0]_net_1 ));
    OR3C \state_RNO_7[0]  (.A(sig_prev), .B(sig_old_i_0), .C(
        \state[0]_net_1 ), .Y(N_270));
    AO1A \state_RNO[0]  (.A(int_enable), .B(\state_ns_0_a2_9[0] ), .C(
        N_26), .Y(\state_ns[0] ));
    DFN1C0 \avg_count[1]  (.D(I_10), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \avg_count[1]_net_1 ));
    NOR2B \count_RNO_0[15]  (.A(count_31_0), .B(count_c13), .Y(N_94));
    NOR3B \state_RNO_3[0]  (.A(\state_ns_0_a2_6[0] ), .B(
        \state_ns_0_a2_5[0] ), .C(avg_enable), .Y(\state_ns_0_a2_8[0] )
        );
    OR3B \state_RNIT6MP[7]  (.A(sig_prev), .B(sig_old_i_0), .C(
        \state[7]_net_1 ), .Y(\state_ns_i_0_0[2] ));
    DFN1E1C0 \count[4]  (.D(count_n4), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[4]_net_1 ));
    DFN1E1C0 \count[12]  (.D(count_n12), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[12]_net_1 ));
    NOR2A \state_RNO[1]  (.A(\state_RNIL4T11[4]_net_1 ), .B(
        next_state15_li), .Y(\state_ns[1] ));
    DFN1E1C0 \count[7]  (.D(count_n7), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[7]_net_1 ));
    
endmodule


module sig_gen_0(
       primary_12_c,
       n_rst_c,
       clk_c,
       sig_old_i_0,
       sig_prev
    );
input  primary_12_c;
input  n_rst_c;
input  clk_c;
output sig_old_i_0;
output sig_prev;

    wire sig_prev_i, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(clk_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev_inst_1 (.D(primary_12_c), .CLK(clk_c), .CLR(
        n_rst_c), .Q(sig_prev));
    INV sig_old_RNO (.A(sig_prev), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module pid_sum_13s_4(
       integral_i,
       integral,
       sr_new,
       sr_new_0_0,
       derivative_0,
       sr_new_1_0,
       integral_0_0,
       integral_1_0,
       sum_39,
       sum_14,
       sum_19,
       sum_20,
       sum_22,
       sum_13,
       sum_18,
       sum_17,
       sum_23,
       sum_21,
       sum_16,
       sum_15,
       sum_12,
       sum_11,
       sum_6,
       sum_10,
       sum_9,
       sum_5,
       sum_8,
       sum_7,
       sum_4,
       sum_2_d0,
       sum_1_d0,
       sum_0_d0,
       sum_3,
       sum_0_0,
       sum_1_0,
       sum_2_0,
       sum_enable,
       sum_rdy,
       n_rst_c,
       clk_c
    );
input  [25:24] integral_i;
input  [25:6] integral;
input  [12:0] sr_new;
input  sr_new_0_0;
input  derivative_0;
input  sr_new_1_0;
input  integral_0_0;
input  integral_1_0;
output sum_39;
output sum_14;
output sum_19;
output sum_20;
output sum_22;
output sum_13;
output sum_18;
output sum_17;
output sum_23;
output sum_21;
output sum_16;
output sum_15;
output sum_12;
output sum_11;
output sum_6;
output sum_10;
output sum_9;
output sum_5;
output sum_8;
output sum_7;
output sum_4;
output sum_2_d0;
output sum_1_d0;
output sum_0_d0;
output sum_3;
output sum_0_0;
output sum_1_0;
output sum_2_0;
input  sum_enable;
output sum_rdy;
input  n_rst_c;
input  clk_c;

    wire \next_sum[39] , \state_RNII1EM[6]_net_1 , \state_0[1]_net_1 , 
        \state_RNIAMDD[0]_net_1 , \state_2[2]_net_1 , 
        \state_1[2]_net_1 , \state_0[2]_net_1 , \state_0[3]_net_1 , 
        \state[6]_net_1 , \un1_next_sum_1_iv_0[26] , 
        next_sum_1_sqmuxa_2, next_sum_1_sqmuxa_1, next_sum_1_sqmuxa, 
        N_416_0, N_12, N_10, \DWACT_FINC_E[0] , N_5, \DWACT_FINC_E[4] , 
        N_2, \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , N_25, N_23, 
        \DWACT_FINC_E_0[0] , N_18, \DWACT_FINC_E_0[4] , N_15, 
        \DWACT_FINC_E_0[7] , \DWACT_FINC_E_0[6] , 
        ADD_40x40_fast_I448_Y_0, \sumreg[30]_net_1 , 
        \un1_next_sum_1_iv[26] , ADD_40x40_fast_I447_Y_0, 
        \sumreg[29]_net_1 , ADD_40x40_fast_I456_Y_0, 
        \sumreg[38]_net_1 , ADD_40x40_fast_I449_Y_0, 
        \sumreg[31]_net_1 , ADD_40x40_fast_I453_Y_0, 
        \sumreg[35]_net_1 , ADD_40x40_fast_I454_Y_0, 
        \sumreg[36]_net_1 , ADD_40x40_fast_I455_Y_0, 
        \sumreg[37]_net_1 , ADD_40x40_fast_I452_Y_0, 
        \sumreg[34]_net_1 , ADD_40x40_fast_I451_Y_0, 
        \sumreg[33]_net_1 , ADD_40x40_fast_I347_Y_0, N787, N772, N771, 
        ADD_40x40_fast_I457_Y_0, ADD_40x40_fast_I446_Y_0, 
        \sumreg[28]_net_1 , ADD_40x40_fast_I450_Y_0, 
        \sumreg[32]_net_1 , ADD_40x40_fast_I348_Y_0, N789, N774, N773, 
        ADD_40x40_fast_I379_Y_4, N840, N871, ADD_40x40_fast_I379_Y_3, 
        N756, ADD_40x40_fast_I379_Y_2, N596, ADD_40x40_fast_I379_Y_0, 
        N681, ADD_40x40_fast_I346_Y_0, N785, N770, N769, 
        ADD_40x40_fast_I382_Y_1, N762, N777, ADD_40x40_fast_I382_Y_0, 
        I194_un1_Y, N687, ADD_40x40_fast_I381_Y_2, N760, N775, 
        ADD_40x40_fast_I381_Y_1, N600, N685, ADD_40x40_fast_I445_Y_0, 
        \sumreg[27]_net_1 , ADD_40x40_fast_I380_Y_2, N758, 
        ADD_40x40_fast_I380_Y_1, I122_un1_Y, N594, N683, 
        ADD_40x40_fast_I432_Y_0, \un1_next_sum_iv_1[14] , 
        \un1_next_sum_iv_2[14] , ADD_40x40_fast_I437_Y_0, 
        \un1_next_sum[19] , ADD_40x40_fast_I438_Y_0, 
        \un1_next_sum[20] , ADD_40x40_fast_I347_un1_Y_0, N788, 
        ADD_40x40_fast_I384_Y_1, N766, N781, ADD_40x40_fast_I384_Y_0, 
        N691, N684, ADD_40x40_fast_I383_Y_1, N764, N779, 
        ADD_40x40_fast_I383_Y_0, N608, N612, ADD_40x40_fast_I443_Y_0, 
        \ireg_m[25] , \un1_next_sum_0_iv_1[25] , \sumreg[25]_net_1 , 
        ADD_40x40_fast_I444_Y_0, \sumreg[26]_net_1 , 
        ADD_40x40_fast_I440_Y_0, \un1_next_sum_2[4] , 
        \un1_next_sum_iv_0[22] , ADD_40x40_fast_I378_Y_4, 
        ADD_40x40_fast_I378_un1_Y_0, N838, ADD_40x40_fast_I378_Y_3, 
        N754, ADD_40x40_fast_I378_Y_2, I118_un1_Y, 
        ADD_40x40_fast_I378_Y_0, ADD_40x40_fast_I431_Y_0, 
        \un1_next_sum_iv_1[13] , \un1_next_sum_iv_2[13] , 
        ADD_40x40_fast_I349_Y_0, I288_un1_Y, ADD_40x40_fast_I385_Y_1, 
        I208_un1_Y, I280_un1_Y, ADD_40x40_fast_I436_Y_0, 
        \un1_next_sum_iv_1[18] , \un1_next_sum_iv_2[18] , 
        ADD_40x40_fast_I435_Y_0, \un1_next_sum_iv_1[17] , 
        \un1_next_sum_iv_2[17] , ADD_40x40_fast_I442_Y_0, 
        \sumreg[24]_net_1 , \un1_next_sum[24] , 
        ADD_40x40_fast_I348_un1_Y_0, N790, ADD_40x40_fast_I441_Y_0, 
        \un1_next_sum[23] , ADD_40x40_fast_I439_Y_0, 
        \un1_next_sum[21] , ADD_40x40_fast_I434_Y_0, 
        \un1_next_sum_iv_1[16] , \un1_next_sum_iv_2[16] , 
        ADD_40x40_fast_I433_Y_0, \un1_next_sum_iv_1[15] , 
        \un1_next_sum_iv_2[15] , ADD_40x40_fast_I346_un1_Y_0, N786, 
        ADD_40x40_fast_I351_Y_0, N795, N780, ADD_40x40_fast_I352_Y_0, 
        N797, N782, ADD_40x40_fast_I430_Y_0, \un1_next_sum_iv_1[12] , 
        \un1_next_sum_iv_2[12] , ADD_40x40_fast_I349_un1_Y_0, N792, 
        N776, ADD_40x40_fast_I353_Y_0, N799, N784, N783, 
        ADD_40x40_fast_I379_un1_Y_0, N804, ADD_40x40_fast_I429_Y_0, 
        \un1_next_sum[11] , ADD_40x40_fast_I424_Y_0, \un1_next_sum[6] , 
        ADD_40x40_fast_I428_Y_0, \un1_next_sum_iv_1[10] , 
        \un1_next_sum_iv_2[10] , ADD_40x40_fast_I427_Y_0, 
        \un1_next_sum[9] , ADD_40x40_fast_I382_un1_Y_0, N743, N878, 
        N802, N817, ADD_40x40_fast_I351_un1_Y_0, N796, 
        ADD_40x40_fast_I352_un1_Y_0, N798, ADD_40x40_fast_I423_Y_0, 
        \un1_next_sum[5] , ADD_40x40_fast_I426_Y_0, 
        \un1_next_sum_iv_1[8] , \un1_next_sum_iv_2[8] , 
        ADD_40x40_fast_I353_un1_Y_0, N800, ADD_40x40_fast_I425_Y_0, 
        \un1_next_sum[7] , ADD_40x40_fast_I383_un1_Y_0, N812, N745, 
        ADD_40x40_fast_I422_Y_0, \un1_next_sum_iv_0[4] , 
        ADD_40x40_fast_I420_Y_0, \un1_next_sum[0] , 
        ADD_40x40_fast_I419_Y_0, ADD_40x40_fast_I257_Y_1, 
        ADD_40x40_fast_I257_Y_0, N661, N472, ADD_40x40_fast_I201_Y_0, 
        N601, N597, ADD_40x40_fast_I197_Y_1, ADD_40x40_fast_I197_Y_0, 
        ADD_40x40_fast_I187_Y_0, ADD_22x22_fast_I126_Y_1, N371, N378, 
        ADD_22x22_fast_I126_Y_0, N335, N332, N331, 
        ADD_22x22_fast_I142_Y_0_1, ADD_22x22_fast_I142_Y_0_a3_0, N329, 
        ADD_22x22_fast_I142_Y_0_0, \i_adj[18]_net_1 , 
        \i_adj[20]_net_1 , N_14_1, ADD_22x22_fast_I172_Y_0, 
        \i_adj[14]_net_1 , \i_adj[12]_net_1 , 
        ADD_22x22_fast_I126_un1_Y_0, N379, 
        ADD_22x22_fast_I142_Y_0_a3_1, N330, ADD_40x40_fast_I418_Y_0, 
        ADD_22x22_fast_I177_Y_0, \i_adj[19]_net_1 , \i_adj[17]_net_1 , 
        ADD_22x22_fast_I178_Y_0, ADD_40x40_fast_I421_Y_0, 
        ADD_22x22_fast_I130_Y_0, N386, ADD_22x22_fast_I142_Y_0_o3_0_0, 
        N337, N334, N333, ADD_22x22_fast_I143_Y_3, 
        ADD_22x22_fast_I143_un1_Y_0, N423, ADD_22x22_fast_I143_Y_2, 
        N367, N374, ADD_22x22_fast_I143_Y_1, N328, 
        ADD_22x22_fast_I143_Y_0, N314, ADD_22x22_fast_I144_Y_2, 
        ADD_22x22_fast_I144_un1_Y_0, N425, ADD_22x22_fast_I144_Y_1, 
        N369, N376, ADD_22x22_fast_I144_Y_0, \un1_next_sum_iv_0[19] , 
        \ireg[19]_net_1 , \un1_next_sum_iv_0[20] , \ireg[20]_net_1 , 
        \un1_next_sum_iv_0[24] , \ireg[24]_net_1 , 
        \un1_next_sum_iv_0[23] , \ireg[23]_net_1 , 
        \un1_next_sum_iv_0[5] , \ireg[5]_net_1 , \ireg[4]_net_1 , 
        \ireg[22]_net_1 , \un1_next_sum_iv_0[21] , \ireg[21]_net_1 , 
        ADD_22x22_fast_I128_Y_0, N382, N375, ADD_22x22_fast_I170_Y_0, 
        \i_adj[10]_net_1 , ADD_22x22_fast_I169_Y_0, \i_adj[11]_net_1 , 
        \i_adj[9]_net_1 , \un24_next_sum_m[12] , next_sum_0_sqmuxa_1, 
        \un3_next_sum_m[12] , \ireg[12]_net_1 , \preg_m[12] , 
        \un24_next_sum_m[18] , \un3_next_sum_m[18] , \ireg[18]_net_1 , 
        \preg_m[18] , \un24_next_sum_m[17] , \un3_next_sum_m[17] , 
        \ireg[17]_net_1 , \preg_m[17] , \un1_next_sum_iv_2[6] , 
        \un3_next_sum_m[6] , \un1_next_sum_iv_0[6] , 
        \un1_next_sum_iv_1[6] , \preg[6]_net_1 , \ireg_m[6] , 
        \un24_next_sum_m[6] , \un24_next_sum_m[13] , 
        \un3_next_sum_m[13] , \preg[13]_net_1 , \ireg_m[13] , 
        \un24_next_sum_m[14] , \un3_next_sum_m[14] , \ireg[14]_net_1 , 
        \preg_m[14] , \un24_next_sum_m[8] , \un3_next_sum_m[8] , 
        \preg[8]_net_1 , \ireg_m[8] , \un24_next_sum_m[10] , 
        \un3_next_sum_m[10] , \preg[10]_net_1 , \ireg_m[10] , 
        \un1_next_sum_iv_2[9] , \un3_next_sum_m[9] , 
        \un1_next_sum_iv_0[9] , \un1_next_sum_iv_1[9] , 
        \preg[9]_net_1 , \ireg_m[9] , \un24_next_sum_m[9] , 
        \un1_next_sum_iv_2[11] , \un24_next_sum_m[11] , 
        \un3_next_sum_m[11] , \un1_next_sum_iv_1[11] , 
        \ireg[11]_net_1 , \preg_m[11] , \un24_next_sum_m[16] , 
        \un3_next_sum_m[16] , \ireg[16]_net_1 , \preg_m[16] , 
        \un24_next_sum_m[15] , \un3_next_sum_m[15] , \ireg[15]_net_1 , 
        \preg_m[15] , \un1_next_sum_iv_2[7] , \un24_next_sum_m[7] , 
        \un3_next_sum_m[7] , \un1_next_sum_iv_1[7] , \preg[7]_net_1 , 
        \ireg_m[7] , next_sum_0_sqmuxa_2, 
        ADD_22x22_fast_I142_Y_0_a3_3_0, N338, ADD_m8_i_1, 
        ADD_m8_i_a4_0_1, N_232, \un3_next_sum_m[25] , 
        ADD_22x22_fast_I129_Y_0, N384, N377, ADD_22x22_fast_I166_Y_0, 
        \i_adj[8]_net_1 , \i_adj[6]_net_1 , 
        ADD_22x22_fast_I128_un1_Y_0, N383, ADD_22x22_fast_I131_Y_0, 
        N345, N342, N341, ADD_22x22_fast_I165_Y_0, \i_adj[7]_net_1 , 
        \i_adj[5]_net_1 , ADD_22x22_fast_I129_un1_Y_0, N385, N266, 
        N359, ADD_22x22_fast_I163_Y_0, \i_adj[3]_net_1 , 
        ADD_22x22_fast_I131_un1_Y_0, N389, N381, N_9, 
        ADD_22x22_fast_I85_Y_0, \i_adj[4]_net_1 , \i_adj[2]_net_1 , 
        N270, ADD_m8_i_o4_1, ADD_m8_i_a4_3, I131_un1_Y, N396, N513, 
        I106_un1_Y, N393, N354, \next_ireg_3[17] , \i_adj[13]_net_1 , 
        \next_ireg_3[11] , N531, \next_ireg_3[16] , N422, I132_un1_Y, 
        \next_ireg_3[14] , N522, \next_ireg_3[7] , \i_adj[1]_net_1 , 
        N682, N1055, N1103, I380_un1_Y, N821, N874, N842, N1025, 
        I334_un1_Y, I383_un1_Y, N848, N1031, I340_un1_Y, N1023, N819, 
        N1040, N1088, N1027, I381_un1_Y, I336_un1_Y, N876, N823, N844, 
        N686, N498, \next_ireg_3[22] , \i_adj[16]_net_1 , 
        \state[5]_net_1 , \state[4]_net_1 , N1037, N1085, N1043, N1091, 
        I382_un1_Y, N778, N1029, I338_un1_Y, \next_ireg_3[25] , 
        \i_adj[21]_net_1 , N492, \next_ireg_3[8] , \next_ireg_3[9] , 
        \next_ireg_3[10] , N394, \next_ireg_3[13] , N525, 
        \next_ireg_3[15] , N424, I133_un1_Y, \next_ireg_3[19] , 
        \i_adj[15]_net_1 , N507, \next_ireg_3[20] , N504, 
        \next_ireg_3[21] , N_11, \next_ireg_3[23] , I124_un1_Y, 
        \next_ireg_3[24] , I122_un1_Y_0, \next_ireg_3[18] , I130_un1_Y, 
        \next_ireg_3[12] , N528, \un1_sumreg[12] , N1094, 
        next_sum_0_sqmuxa, N1035, I385_un1_Y, I344_un1_Y, N884, N852, 
        N1033, I384_un1_Y, I342_un1_Y, N882, N666, N850, N1058, N1106, 
        N1052, N1100, N1049, I290_un1_Y, I350_un1_Y, N794, N1097, 
        N1046, N595, N599, N591, N680, N387, N1021, N869, 
        \state[1]_net_1 , N740, N659, \inf_abs1_5[0] , \inf_abs1_5[2] , 
        \inf_abs1_a_2[2] , \inf_abs1_5[3] , \inf_abs1_a_2[3] , 
        \inf_abs1_5[4] , \inf_abs1_a_2[4] , \inf_abs1_5[5] , 
        \inf_abs1_a_2[5] , \inf_abs1_5[7] , \inf_abs1_a_2[7] , 
        \inf_abs1_5[9] , \inf_abs1_a_2[9] , \inf_abs1_5[10] , 
        \inf_abs1_a_2[10] , \inf_abs1_5[11] , \inf_abs1_a_2[11] , 
        \inf_abs2_5[0] , \inf_abs2_5[2] , \inf_abs2_a_0[2] , 
        \inf_abs2_5[14] , \inf_abs2_a_0[14] , \state[2]_net_1 , 
        \inf_abs2_5[12] , \inf_abs2_a_0[12] , \next_sum[1] , 
        \next_sum[2] , \next_sum[5] , \next_sum[6] , \next_sum[8] , 
        \next_sum[12] , \next_sum[13] , \next_sum[14] , \next_sum[15] , 
        \next_sum[16] , N1082, \next_sum[17] , N1079, \next_sum[18] , 
        N1076, \next_sum[21] , N1067, \next_sum[22] , N1064, 
        \next_sum[23] , N1061, \next_sum[24] , \next_sum[26] , 
        \next_sum[27] , \next_sum[28] , \next_sum[32] , \next_sum[33] , 
        N282, N284, N288, N347, N287, N351, N278, N281, N352, N279, 
        N344, N343, N348, N390, N355, N391, N356, I114_un1_Y, N350, 
        N340, N336, N305, N308, N311, N312, N309, N392, 
        \next_ireg_3[6] , \i_adj[0]_net_1 , N388, N349, N725, N648, 
        N645, N644, N726, N649, I116_un1_Y, N664, I216_un1_Y, N701, 
        N694, N693, N702, N709, N710, I232_un1_Y, N717, N791, N641, 
        N637, I240_un1_Y, N807, N733, I252_un1_Y, N653, N737, N811, 
        N729, N738, I256_un1_Y, N741, N734, I359_un1_Y, I308_un1_Y, 
        I361_un1_Y, N883, N490, N493, N713, N636, N633, N632, N519, 
        N523, N522_0, N520, N621, N538, N541, N706, N625, N629, N529, 
        N526, N657, N660, N628, N525_0, N528_0, N624, N620, N537, N540, 
        N613, N616, N652, N489, N492_0, N499, N496, N486, N487, N507_0, 
        N508, N514, N642, N504_0, N643, N505, N650, N495, N651, N654, 
        N655, N716, N639, N635, I166_un1_Y, N719, N638, N720, N723, 
        N646, N724, N647, N727, N728, N731, N732, N735, N658, N736, 
        N739, N662, N704, N712, N793, N711, N801, N806, N809, N810, 
        I254_un1_Y, N814, N877, N631, N634, N630, N513_0, N516, N517, 
        N534, N543, N544, N618, N619, N607, N603, N610, N606, N688, 
        N611, N614, N692, N615, N695, N697, N617, N623, N627, N705, 
        N707, N626, N708, N715, N696, N699, N700, N703, N805, N808, 
        I300_un1_Y, N803, I302_un1_Y, N873, I310_un1_Y, I320_un1_Y, 
        I354_un1_Y, I355_un1_Y, I360_un1_Y, \inf_abs2_5[6] , 
        \inf_abs2_a_0[6] , \inf_abs2_5[15] , \inf_abs2_a_0[15] , 
        \inf_abs2_5[16] , \inf_abs2_a_0[16] , \inf_abs2_5[18] , 
        \inf_abs2_a_0[18] , \inf_abs2_5[19] , \inf_abs2_a_0[19] , 
        \inf_abs2_5[20] , \inf_abs2_a_0[20] , \inf_abs2_5[21] , 
        \inf_abs2_a_0[21] , \state[3]_net_1 , \ireg[6]_net_1 , 
        \ireg[7]_net_1 , \ireg[8]_net_1 , \ireg[9]_net_1 , 
        \ireg[10]_net_1 , \preg[12]_net_1 , \ireg[13]_net_1 , 
        \preg[14]_net_1 , \preg[15]_net_1 , \preg[16]_net_1 , 
        \preg[17]_net_1 , \preg[18]_net_1 , \ireg[25]_net_1 , N339, 
        N602, \next_sum[35] , N481, N480, N484, N483, N656, 
        \next_sum[29] , \next_sum[4] , \next_sum[3] , I244_un1_Y, N722, 
        N875, N721, N714, I321_un1_Y, I312_un1_Y, \next_sum[31] , 
        N_228, \inf_abs1_5[1] , \inf_abs1_a_2[1] , N471, \next_sum[0] , 
        \state_ns[0] , \inf_abs1_5[12] , \inf_abs1_a_2[12] , 
        \inf_abs1_5[6] , \inf_abs1_a_2[6] , \inf_abs1_5[8] , 
        \inf_abs1_a_2[8] , N502, N501, N498_0, \next_sum[10] , 
        \preg[11]_net_1 , N1073, I358_un1_Y, I298_un1_Y, I168_un1_Y, 
        N640, N622, N511, N510, \next_sum[19] , \next_sum[11] , 
        \next_sum[9] , \next_sum[7] , N1070, N532, N531_0, 
        \next_sum[20] , \next_sum[36] , N604, N605, N609, 
        \next_sum[30] , \next_sum[38] , N698, N690, I212_un1_Y, N547, 
        N546, \next_sum[37] , \next_sum[34] , \next_sum[25] , 
        \inf_abs2_5[17] , \inf_abs2_a_0[17] , \inf_abs2_5[11] , 
        \inf_abs2_a_0[11] , \inf_abs2_5[8] , \inf_abs2_a_0[8] , 
        \inf_abs2_5[5] , \inf_abs2_a_0[5] , \inf_abs2_5[7] , 
        \inf_abs2_a_0[7] , \inf_abs2_5[4] , \inf_abs2_a_0[4] , 
        \inf_abs2_5[13] , \inf_abs2_a_0[13] , \inf_abs2_5[10] , 
        \inf_abs2_a_0[10] , \inf_abs2_5[9] , \inf_abs2_a_0[9] , 
        \inf_abs2_5[3] , \inf_abs2_a_0[3] , \inf_abs2_5[1] , 
        \inf_abs2_a_0[1] , N297, N291, N290, N353, N275, N357, N269, 
        I115_un1_Y, I54_un1_Y, N346, N303, N299, N302, N306, N296, 
        N293, N294, N276, N272, \p_adj[0]_net_1 , \p_adj[1]_net_1 , 
        \p_adj[2]_net_1 , \p_adj[3]_net_1 , \p_adj[4]_net_1 , 
        \p_adj[5]_net_1 , \p_adj[6]_net_1 , \p_adj[7]_net_1 , 
        \p_adj[8]_net_1 , \p_adj[9]_net_1 , \p_adj[10]_net_1 , 
        \p_adj[11]_net_1 , \p_adj[12]_net_1 , N_6, \DWACT_FINC_E[28] , 
        \DWACT_FINC_E[13] , \DWACT_FINC_E[15] , N_7, 
        \DWACT_FINC_E[14] , N_8, \DWACT_FINC_E[9] , \DWACT_FINC_E[12] , 
        N_9_0, \DWACT_FINC_E[10] , \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[5] , N_10_0, \DWACT_FINC_E[11] , N_11_0, N_12_0, 
        N_13, \DWACT_FINC_E[8] , N_14, N_16, N_17, \DWACT_FINC_E[3] , 
        N_19, N_20, N_21, \DWACT_FINC_E[1] , N_22, N_24, N_3, 
        \DWACT_FINC_E_0[2] , \DWACT_FINC_E_0[5] , N_4, 
        \DWACT_FINC_E_0[3] , N_6_0, N_7_0, N_8_0, \DWACT_FINC_E_0[1] , 
        N_9_1, N_11_1, GND, VCC;
    
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I312_un1_Y (.A(N733), .B(
        I256_un1_Y), .C(N800), .Y(I312_un1_Y));
    DFN1E1C0 \sumreg[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(sum_39));
    NOR3B \preg_RNIJKQK[7]  (.A(sr_new_0_0), .B(\state[5]_net_1 ), .C(
        \preg[7]_net_1 ), .Y(\un24_next_sum_m[7] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I77_Y (.A(N532), .B(N529), .Y(
        N627));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_o3_0 (.A(
        ADD_22x22_fast_I142_Y_0_a3_3_0), .B(N513), .C(
        ADD_22x22_fast_I142_Y_0_o3_0_0), .Y(N_11));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I19_G0N (.A(\un1_next_sum[19] )
        , .B(sum_19), .Y(N528_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I14_P0N (.A(
        \un1_next_sum_iv_1[14] ), .B(\un1_next_sum_iv_2[14] ), .C(
        sum_14), .Y(N514));
    OR3 \ireg_RNIN85P1[12]  (.A(\un24_next_sum_m[12] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[12] ), .Y(
        \un1_next_sum_iv_2[12] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I46_Y (.A(\sumreg[34]_net_1 ), 
        .B(\sumreg[35]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N596)
        );
    XA1B \sumreg_RNO[10]  (.A(N1100), .B(ADD_40x40_fast_I428_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[10] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I118_un1_Y (.A(N591), .B(N594), 
        .Y(I118_un1_Y));
    MX2 \p_adj_RNO[2]  (.A(sr_new[2]), .B(\inf_abs1_a_2[2] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[2] ));
    AO1 \ireg_RNIDJU91[12]  (.A(\ireg[12]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[12] ), .Y(
        \un1_next_sum_iv_1[12] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I336_un1_Y (.A(N844), .B(N875), 
        .Y(I336_un1_Y));
    XA1B \sumreg_RNO[11]  (.A(N1097), .B(ADD_40x40_fast_I429_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[11] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_0 (.A(N333), .B(N330), .C(
        N329), .Y(ADD_22x22_fast_I144_Y_0));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I241_Y (.A(N641), .B(N637), .C(
        N726), .Y(N800));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I114_Y (.A(N471), .B(
        \un1_next_sum[0] ), .C(sum_1_d0), .Y(N664));
    DFN1E1C0 \i_adj[19]  (.D(\inf_abs2_5[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[19]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I113_Y (.A(N389), .B(N396), .C(
        N388), .Y(N525));
    DFN1E1C0 \sumreg[23]  (.D(\next_sum[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(sum_23));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I290_un1_Y (.A(N793), .B(N778), 
        .Y(I290_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I128_un1_Y_0 (.A(N383), .B(N375)
        , .Y(ADD_22x22_fast_I128_un1_Y_0));
    NOR3B inf_abs1_a_2_I_19 (.A(\DWACT_FINC_E_0[2] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[6]), .Y(N_7_0));
    OA1 next_ireg_3_0_ADD_22x22_fast_I33_Y (.A(\i_adj[11]_net_1 ), .B(
        \i_adj[13]_net_1 ), .C(N303), .Y(N338));
    NOR2B \preg_RNILLAM[17]  (.A(\preg[17]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[17] ));
    AND3 inf_abs2_a_0_I_30 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E_0[6] ));
    MX2 \i_adj_RNO[5]  (.A(integral[11]), .B(\inf_abs2_a_0[5] ), .S(
        integral_0_0), .Y(\inf_abs2_5[5] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I304_Y (.A(N807), .B(N792), .C(
        N791), .Y(N875));
    DFN1E1C0 \sumreg[38]  (.D(\next_sum[38] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[38]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I126_un1_Y_0 (.A(N371), .B(N379)
        , .Y(ADD_22x22_fast_I126_un1_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I361_Y (.A(I361_un1_Y), .B(N883), 
        .Y(N1082));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I201_Y_0 (.A(N601), .B(N597), 
        .Y(ADD_40x40_fast_I201_Y_0));
    DFN1E1C0 \sumreg[5]  (.D(\next_sum[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_5));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I248_Y (.A(N733), .B(N726), .C(
        N725), .Y(N807));
    DFN1E1C0 \sumreg[20]  (.D(\next_sum[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(sum_20));
    AO1 next_ireg_3_0_ADD_22x22_fast_I128_Y (.A(
        ADD_22x22_fast_I128_un1_Y_0), .B(N528), .C(
        ADD_22x22_fast_I128_Y_0), .Y(N504));
    OR2 \preg_RNISQKN2[9]  (.A(\un1_next_sum_iv_2[9] ), .B(
        \un1_next_sum_iv_1[9] ), .Y(\un1_next_sum[9] ));
    NOR2 inf_abs2_a_0_I_57 (.A(integral[24]), .B(integral[25]), .Y(
        \DWACT_FINC_E[14] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I347_Y_0 (.A(N787), .B(N772), .C(
        N771), .Y(ADD_40x40_fast_I347_Y_0));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I52_Y (.A(\sumreg[32]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N602)
        );
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I199_Y (.A(N595), .B(N599), .C(
        N684), .Y(N758));
    DFN1E1C0 \sumreg[13]  (.D(\next_sum[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_13));
    XA1 \ireg_RNISPNG[21]  (.A(integral_1_0), .B(\ireg[21]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[21] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I354_Y (.A(I354_un1_Y), .B(N869), 
        .Y(N1061));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I214_Y (.A(N699), .B(N692), .C(
        N691), .Y(N773));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I353_un1_Y_0 (.A(N800), .B(
        N784), .Y(ADD_40x40_fast_I353_un1_Y_0));
    DFN1E1C0 \i_adj[2]  (.D(\inf_abs2_5[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[2]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I225_Y (.A(N702), .B(N710), .Y(
        N784));
    NOR3A inf_abs1_a_2_I_13 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .C(
        sr_new[4]), .Y(N_9_1));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I436_Y_0 (.A(
        \un1_next_sum_iv_1[18] ), .B(\un1_next_sum_iv_2[18] ), .C(
        sum_18), .Y(ADD_40x40_fast_I436_Y_0));
    DFN1E1C0 \sumreg[27]  (.D(\next_sum[27] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[27]_net_1 ));
    DFN1E1C0 \sumreg[10]  (.D(\next_sum[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_10));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I381_Y_2 (.A(N760), .B(N775), .C(
        ADD_40x40_fast_I381_Y_1), .Y(ADD_40x40_fast_I381_Y_2));
    XA1 \ireg_RNIRONG[20]  (.A(integral_1_0), .B(\ireg[20]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[20] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I15_P0N (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(N312));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I444_Y_0 (.A(
        \sumreg[26]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I444_Y_0));
    XA1B \sumreg_RNO[22]  (.A(N1064), .B(ADD_40x40_fast_I440_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[22] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I171_Y (.A(N647), .B(N643), .Y(
        N724));
    AX1B un1_sumreg_0_0_ADD_40x40_fast_I443_Y_0 (.A(\ireg_m[25] ), .B(
        \un1_next_sum_0_iv_1[25] ), .C(\sumreg[25]_net_1 ), .Y(
        ADD_40x40_fast_I443_Y_0));
    AND2 inf_abs2_a_0_I_44 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E[9] ), .Y(\DWACT_FINC_E[10] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I18_P0N (.A(
        \un1_next_sum_iv_1[18] ), .B(\un1_next_sum_iv_2[18] ), .C(
        sum_18), .Y(N526));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I166_Y (.A(I166_un1_Y), .B(N638), 
        .Y(N719));
    OR2 \preg_RNIKIKN2[7]  (.A(\un1_next_sum_iv_2[7] ), .B(
        \un1_next_sum_iv_1[7] ), .Y(\un1_next_sum[7] ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_0_0 (.A(
        \i_adj[18]_net_1 ), .B(\i_adj[20]_net_1 ), .C(N_9), .Y(
        ADD_22x22_fast_I142_Y_0_a3_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I10_P0N (.A(\i_adj[12]_net_1 ), 
        .B(\i_adj[10]_net_1 ), .Y(N297));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I168_Y (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[8]_net_1 ), .C(N522), .Y(\next_ireg_3[14] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I384_Y_1 (.A(N766), .B(N781), .C(
        ADD_40x40_fast_I384_Y_0), .Y(ADD_40x40_fast_I384_Y_1));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I10_G0N (.A(
        \un1_next_sum_iv_1[10] ), .B(\un1_next_sum_iv_2[10] ), .C(
        sum_10), .Y(N501));
    XNOR2 inf_abs1_a_2_I_28 (.A(sr_new[10]), .B(N_4), .Y(
        \inf_abs1_a_2[10] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I18_G0N (.A(
        \un1_next_sum_iv_1[18] ), .B(\un1_next_sum_iv_2[18] ), .C(
        sum_18), .Y(N525_0));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I338_un1_Y (.A(N778), .B(N762), 
        .C(N877), .Y(I338_un1_Y));
    DFN1E1C0 \p_adj[4]  (.D(\inf_abs1_5[4] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[4]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_2 (.A(
        ADD_22x22_fast_I144_un1_Y_0), .B(N425), .C(
        ADD_22x22_fast_I144_Y_1), .Y(ADD_22x22_fast_I144_Y_2));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I358_Y (.A(I358_un1_Y), .B(N877), 
        .Y(N1073));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I7_G0N (.A(\i_adj[9]_net_1 ), 
        .B(\i_adj[7]_net_1 ), .Y(N287));
    XNOR2 inf_abs2_a_0_I_20 (.A(integral[13]), .B(N_20), .Y(
        \inf_abs2_a_0[7] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I424_Y_0 (.A(sum_6), .B(
        \un1_next_sum[6] ), .Y(ADD_40x40_fast_I424_Y_0));
    DFN1E1C0 \sumreg[17]  (.D(\next_sum[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_17));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I257_Y_1 (.A(
        ADD_40x40_fast_I257_Y_0), .B(N661), .Y(ADD_40x40_fast_I257_Y_1)
        );
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I321_Y (.A(N733), .B(I256_un1_Y), 
        .C(I321_un1_Y), .Y(N1106));
    DFN1C0 \state[6]  (.D(\state_1[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[6]_net_1 ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I423_Y_0 (.A(sum_5), .B(
        \un1_next_sum[5] ), .Y(ADD_40x40_fast_I423_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y (.A(
        ADD_22x22_fast_I126_un1_Y_0), .B(N522), .C(
        ADD_22x22_fast_I126_Y_1), .Y(N498));
    AND3 inf_abs1_a_2_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[5] ), .Y(
        \DWACT_FINC_E[6] ));
    DFN1E1C0 \sumreg[35]  (.D(\next_sum[35] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[35]_net_1 ));
    MX2 \i_adj_RNO[13]  (.A(integral[19]), .B(\inf_abs2_a_0[13] ), .S(
        integral_0_0), .Y(\inf_abs2_5[13] ));
    DFN1E1C0 \sumreg[4]  (.D(\next_sum[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_4));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I166_Y_0 (.A(\i_adj[8]_net_1 ), 
        .B(\i_adj[6]_net_1 ), .Y(ADD_22x22_fast_I166_Y_0));
    XA1B \sumreg_RNO[38]  (.A(N1023), .B(ADD_40x40_fast_I456_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[38] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I160_Y (.A(N636), .B(N633), .C(
        N632), .Y(N713));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I342_un1_Y (.A(N797), .B(
        I310_un1_Y), .C(N850), .Y(I342_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I207_Y (.A(N684), .B(N692), .Y(
        N766));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I232_Y (.A(I232_un1_Y), .B(N709), 
        .Y(N791));
    NOR2 inf_abs2_a_0_I_6 (.A(integral[6]), .B(integral[7]), .Y(N_25));
    NOR3B inf_abs2_a_0_I_45 (.A(\DWACT_FINC_E[10] ), .B(
        \DWACT_FINC_E_0[6] ), .C(integral[21]), .Y(N_11_0));
    NOR2A \state_RNINQBC_0[5]  (.A(\state[5]_net_1 ), .B(sr_new[12]), 
        .Y(next_sum_1_sqmuxa_2));
    XA1 \ireg_RNIVSNG[24]  (.A(integral_1_0), .B(\ireg[24]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[24] ));
    NOR3 inf_abs1_a_2_I_29 (.A(sr_new[7]), .B(sr_new[6]), .C(sr_new[8])
        , .Y(\DWACT_FINC_E_0[5] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I252_Y (.A(I252_un1_Y), .B(N729), 
        .Y(N811));
    MX2 \p_adj_RNO[1]  (.A(sr_new[1]), .B(\inf_abs1_a_2[1] ), .S(
        sr_new_1_0), .Y(\inf_abs1_5[1] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I382_un1_Y (.A(N778), .B(N762), 
        .C(ADD_40x40_fast_I382_un1_Y_0), .Y(I382_un1_Y));
    NOR3B \preg_RNIGGAM[12]  (.A(\state[5]_net_1 ), .B(
        \preg[12]_net_1 ), .C(sr_new[12]), .Y(\preg_m[12] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I252_un1_Y (.A(N653), .B(N649), 
        .C(N737), .Y(I252_un1_Y));
    AO1 next_ireg_3_0_ADD_22x22_fast_I30_Y (.A(N302), .B(N306), .C(
        N305), .Y(N335));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I124_un1_Y (.A(N377), .B(N369), 
        .C(N424), .Y(I124_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I237_Y (.A(N714), .B(N722), .Y(
        N796));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I12_G0N (.A(\i_adj[12]_net_1 ), 
        .B(\i_adj[14]_net_1 ), .Y(N302));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I11_G0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(N299));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I58_Y (.A(\sumreg[28]_net_1 ), 
        .B(\sumreg[29]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N608)
        );
    OA1 next_ireg_3_0_ADD_22x22_fast_I35_Y (.A(\i_adj[11]_net_1 ), .B(
        \i_adj[13]_net_1 ), .C(N297), .Y(N340));
    DFN1E1C0 \sumreg[7]  (.D(\next_sum[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_7));
    DFN1E1C0 \ireg[12]  (.D(\next_ireg_3[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[12]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I126_Y (.A(N602), .B(I122_un1_Y), 
        .Y(I194_un1_Y));
    NOR2A inf_abs2_a_0_I_11 (.A(\DWACT_FINC_E_0[0] ), .B(integral[9]), 
        .Y(N_23));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I197_Y_1 (.A(
        ADD_40x40_fast_I197_Y_0), .B(N597), .Y(ADD_40x40_fast_I197_Y_1)
        );
    XOR2 next_ireg_3_0_ADD_22x22_fast_I166_Y (.A(
        ADD_22x22_fast_I166_Y_0), .B(N528), .Y(\next_ireg_3[12] ));
    AO1 \preg_RNIJ9R41[6]  (.A(\preg[6]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[6] ), .Y(
        \un1_next_sum_iv_1[6] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I67_Y (.A(N547), .B(N544), .Y(
        N617));
    AO1 next_ireg_3_0_ADD_22x22_fast_I38_Y (.A(N290), .B(N294), .C(
        N293), .Y(N343));
    XNOR2 inf_abs2_a_0_I_46 (.A(integral[22]), .B(N_11_0), .Y(
        \inf_abs2_a_0[16] ));
    XOR2 inf_abs1_a_2_I_5 (.A(sr_new[0]), .B(sr_new[1]), .Y(
        \inf_abs1_a_2[1] ));
    XNOR2 inf_abs1_a_2_I_23 (.A(sr_new[8]), .B(N_6_0), .Y(
        \inf_abs1_a_2[8] ));
    NOR3B \preg_RNIUDN01[10]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), 
        .C(\preg[10]_net_1 ), .Y(\un24_next_sum_m[10] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I308_un1_Y (.A(N811), .B(N796), 
        .Y(I308_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I169_Y (.A(N641), .B(N645), .Y(
        N722));
    DFN1C0 \state[2]  (.D(\state[1]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[2]_net_1 ));
    OR2 \ireg_RNIEKQ41[21]  (.A(\un1_next_sum_iv_0[21] ), .B(
        \un1_next_sum_2[4] ), .Y(\un1_next_sum[21] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I245_Y (.A(N653), .B(N649), .C(
        N722), .Y(N804));
    DFN1E1C0 \i_adj[15]  (.D(\inf_abs2_5[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[15]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I349_Y_0 (.A(N775), .B(
        I288_un1_Y), .Y(ADD_40x40_fast_I349_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I41_Y (.A(N291), .B(N288), .Y(
        N346));
    DFN1E1C0 \i_adj[20]  (.D(\inf_abs2_5[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[20]_net_1 ));
    XNOR2 inf_abs2_a_0_I_37 (.A(integral[19]), .B(N_14), .Y(
        \inf_abs2_a_0[13] ));
    MX2 \i_adj_RNO[12]  (.A(integral[18]), .B(\inf_abs2_a_0[12] ), .S(
        integral_0_0), .Y(\inf_abs2_5[12] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I348_Y_0 (.A(N789), .B(N774), .C(
        N773), .Y(ADD_40x40_fast_I348_Y_0));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I53_Y (.A(\sumreg[32]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N603)
        );
    AO1 next_ireg_3_0_ADD_22x22_fast_I86_Y (.A(N356), .B(N359), .C(
        N355), .Y(N394));
    NOR2B \preg_RNIKKAM[16]  (.A(\preg[16]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[16] ));
    AX1D next_ireg_3_0_ADD_22x22_fast_I170_Y (.A(N422), .B(I132_un1_Y), 
        .C(ADD_22x22_fast_I170_Y_0), .Y(\next_ireg_3[16] ));
    AO1 \preg_RNILBR41[7]  (.A(\preg[7]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[7] ), .Y(
        \un1_next_sum_iv_1[7] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_1 (.A(N369), .B(N376), .C(
        ADD_22x22_fast_I144_Y_0), .Y(ADD_22x22_fast_I144_Y_1));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I4_P0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[4] ), .C(sum_4), .Y(N484));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I213_Y (.A(N690), .B(N698), .Y(
        N772));
    NOR3 \state_RNI1KGU[6]  (.A(sum_rdy), .B(\state[6]_net_1 ), .C(
        \state_0[1]_net_1 ), .Y(N_416_0));
    DFN1E1C0 \p_adj[10]  (.D(\inf_abs1_5[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[10]_net_1 ));
    DFN1E1C0 \p_adj[5]  (.D(\inf_abs1_5[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[5]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I164_Y (.A(N640), .B(N637), .C(
        N636), .Y(N717));
    DFN1E1C0 \sumreg[36]  (.D(\next_sum[36] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[36]_net_1 ));
    NOR3B \preg_RNIKLQK[8]  (.A(sr_new_0_0), .B(\state[5]_net_1 ), .C(
        \preg[8]_net_1 ), .Y(\un24_next_sum_m[8] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I56_Y (.A(\sumreg[29]_net_1 ), 
        .B(\sumreg[30]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N606)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I172_Y (.A(N648), .B(N645), .C(
        N644), .Y(N725));
    NOR2B \p_adj_RNO[12]  (.A(\inf_abs1_a_2[12] ), .B(sr_new[12]), .Y(
        \inf_abs1_5[12] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I300_un1_Y (.A(N803), .B(N788), 
        .Y(I300_un1_Y));
    DFN1E1C0 \p_adj[0]  (.D(\inf_abs1_5[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[0]_net_1 ));
    AND3 inf_abs2_a_0_I_51 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[28] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I354_un1_Y (.A(N786), .B(N802), 
        .C(N817), .Y(I354_un1_Y));
    OR2 \preg_RNI0IKC2[6]  (.A(\un1_next_sum_iv_2[6] ), .B(
        \un1_next_sum_iv_1[6] ), .Y(\un1_next_sum[6] ));
    DFN1E1C0 \sumreg[9]  (.D(\next_sum[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_9));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I181_Y (.A(N657), .B(N653), .Y(
        N734));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I216_Y (.A(I216_un1_Y), .B(N693), 
        .Y(N775));
    NOR3B \preg_RNI1HN01[13]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), 
        .C(\preg[13]_net_1 ), .Y(\un24_next_sum_m[13] ));
    OA1 un1_sumreg_0_0_ADD_m8_i_a4 (.A(N_232), .B(ADD_m8_i_o4_1), .C(
        next_sum_0_sqmuxa), .Y(ADD_m8_i_a4_3));
    NOR3B \ireg_RNISOMG[12]  (.A(integral_1_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[12]_net_1 ), .Y(\un3_next_sum_m[12] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I4_G0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[4] ), .C(sum_4), .Y(N483));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I317_Y (.A(N808), .B(N823), .C(
        N807), .Y(N1094));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I129_Y (.A(N605), .B(N601), .Y(
        N682));
    NOR3B \ireg_RNIGH7M[6]  (.A(\state[3]_net_1 ), .B(\ireg[6]_net_1 ), 
        .C(integral[25]), .Y(\ireg_m[6] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I50_Y (.A(N272), .B(N276), .C(
        N275), .Y(N355));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I144_un1_Y_0 (.A(N377), .B(N369)
        , .C(N266), .Y(ADD_22x22_fast_I144_un1_Y_0));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I34_Y (.A(N296), .B(
        \i_adj[11]_net_1 ), .C(\i_adj[13]_net_1 ), .Y(N339));
    DFN1E1C0 \sumreg[31]  (.D(\next_sum[31] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[31]_net_1 ));
    NOR3B \preg_RNIIJQK[6]  (.A(sr_new_0_0), .B(\state[5]_net_1 ), .C(
        \preg[6]_net_1 ), .Y(\un24_next_sum_m[6] ));
    DFN1E1C0 \sumreg[2]  (.D(\next_sum[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_2_d0));
    DFN1E1C0 \i_adj[7]  (.D(\inf_abs2_5[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[7]_net_1 ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I383_Y (.A(
        ADD_40x40_fast_I383_Y_1), .B(I383_un1_Y), .C(I340_un1_Y), .Y(
        N1031));
    MX2 \i_adj_RNO[8]  (.A(integral[14]), .B(\inf_abs2_a_0[8] ), .S(
        integral_0_0), .Y(\inf_abs2_5[8] ));
    AO1 \ireg_RNILRU91[16]  (.A(\ireg[16]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[16] ), .Y(
        \un1_next_sum_iv_1[16] ));
    AO1 \preg_RNI85171[10]  (.A(\preg[10]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[10] ), .Y(
        \un1_next_sum_iv_1[10] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I9_P0N (.A(\un1_next_sum[9] ), 
        .B(sum_9), .Y(N499));
    NOR3A inf_abs2_a_0_I_27 (.A(\DWACT_FINC_E_0[4] ), .B(integral[14]), 
        .C(integral[15]), .Y(N_17));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I105_Y (.A(N487), .B(N490), .Y(
        N655));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I10_G0N (.A(\i_adj[12]_net_1 ), 
        .B(\i_adj[10]_net_1 ), .Y(N296));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I351_un1_Y_0 (.A(N796), .B(
        N780), .Y(ADD_40x40_fast_I351_un1_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I108_Y (.A(N390), .B(N383), .C(
        N382), .Y(N422));
    MX2 \p_adj_RNO[3]  (.A(sr_new[3]), .B(\inf_abs1_a_2[3] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[3] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I435_Y_0 (.A(
        \un1_next_sum_iv_1[17] ), .B(\un1_next_sum_iv_2[17] ), .C(
        sum_17), .Y(ADD_40x40_fast_I435_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I146_Y (.A(N622), .B(N619), .C(
        N618), .Y(N699));
    AND3 inf_abs2_a_0_I_48 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[11] ), .Y(N_10_0));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I197_Y_0 (.A(\sumreg[36]_net_1 )
        , .B(\sumreg[37]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(
        ADD_40x40_fast_I197_Y_0));
    DFN1E1C0 \preg[16]  (.D(\p_adj[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[16]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I135_Y (.A(N611), .B(N607), .Y(
        N688));
    NOR3B \preg_RNI4KN01[16]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), 
        .C(\preg[16]_net_1 ), .Y(\un24_next_sum_m[16] ));
    DFN1E1C0 \preg[17]  (.D(\p_adj[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[17]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I9_G0N (.A(\i_adj[9]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(N293));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I155_Y (.A(N627), .B(N631), .Y(
        N708));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I122_un1_Y (.A(N375), .B(N367), 
        .C(N422), .Y(I122_un1_Y_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I12_P0N (.A(\i_adj[12]_net_1 ), 
        .B(\i_adj[14]_net_1 ), .Y(N303));
    OR2 next_ireg_3_0_ADD_22x22_fast_I5_P0N (.A(\i_adj[5]_net_1 ), .B(
        \i_adj[7]_net_1 ), .Y(N282));
    DFN1E1C0 \i_adj[8]  (.D(\inf_abs2_5[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[8]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I94_Y (.A(N501), .B(N505), .C(
        N504_0), .Y(N644));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I73_Y (.A(N342), .B(N346), .Y(
        N381));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I174_Y (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .C(N504), .Y(\next_ireg_3[20] ));
    DFN1E1C0 \i_adj[17]  (.D(\inf_abs2_5[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[17]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I140_Y (.A(N616), .B(N613), .C(
        N612), .Y(N693));
    MX2 \i_adj_RNO[3]  (.A(integral[9]), .B(\inf_abs2_a_0[3] ), .S(
        integral_0_0), .Y(\inf_abs2_5[3] ));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I74_Y (.A(N531_0), .B(sum_21), 
        .C(\un1_next_sum[21] ), .Y(N624));
    XNOR2 inf_abs2_a_0_I_49 (.A(integral[23]), .B(N_10_0), .Y(
        \inf_abs2_a_0[17] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I168_un1_Y (.A(N644), .B(N641), 
        .Y(I168_un1_Y));
    XNOR2 inf_abs2_a_0_I_12 (.A(integral[10]), .B(N_23), .Y(
        \inf_abs2_a_0[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I319_Y (.A(N812), .B(N745), .C(
        N811), .Y(N1100));
    XA1B \sumreg_RNO[18]  (.A(N1076), .B(ADD_40x40_fast_I436_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[18] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I383_un1_Y_0 (.A(N796), .B(
        N812), .C(N745), .Y(ADD_40x40_fast_I383_un1_Y_0));
    AO1 \preg_RNIEB171[13]  (.A(\preg[13]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[13] ), .Y(
        \un1_next_sum_iv_1[13] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I306_Y (.A(N809), .B(N794), .C(
        N793), .Y(N877));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I224_Y (.A(N709), .B(N702), .C(
        N701), .Y(N783));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I383_Y_0 (.A(N608), .B(N612), .C(
        N681), .Y(ADD_40x40_fast_I383_Y_0));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I17_G0N (.A(
        \un1_next_sum_iv_1[17] ), .B(\un1_next_sum_iv_2[17] ), .C(
        sum_17), .Y(N522_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I356_Y (.A(N874), .B(N821), .C(
        N873), .Y(N1067));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I239_Y (.A(N716), .B(N724), .Y(
        N798));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I259_Y (.A(N738), .B(N745), .C(
        N737), .Y(N819));
    NOR2B \i_adj_RNO[21]  (.A(\inf_abs2_a_0[21] ), .B(integral[25]), 
        .Y(\inf_abs2_5[21] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I116_un1_Y (.A(N472), .B(
        \un1_next_sum[0] ), .Y(I116_un1_Y));
    DFN1E1C0 \sumreg[6]  (.D(\next_sum[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_6));
    DFN1E1C0 \sumreg[0]  (.D(\next_sum[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_0_d0));
    DFN1E1C0 \preg[15]  (.D(\p_adj[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[15]_net_1 ));
    DFN1E1C0 \i_adj[10]  (.D(\inf_abs2_5[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[10]_net_1 ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I452_Y_0 (.A(
        \sumreg[34]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I452_Y_0));
    DFN1E1C0 \ireg[24]  (.D(\next_ireg_3[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[24]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I271_Y (.A(N758), .B(N774), .Y(
        N842));
    NOR2A \ireg_RNI18LJ_0[25]  (.A(next_sum_1_sqmuxa), .B(
        \ireg[25]_net_1 ), .Y(\un3_next_sum_m[25] ));
    XNOR2 inf_abs2_a_0_I_43 (.A(integral[21]), .B(N_12_0), .Y(
        \inf_abs2_a_0[15] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I69_Y (.A(N342), .B(N338), .Y(
        N377));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I385_Y (.A(I385_un1_Y), .B(
        ADD_40x40_fast_I385_Y_1), .C(I344_un1_Y), .Y(N1035));
    NOR3B \ireg_RNIG9K8[15]  (.A(integral_1_0), .B(\state[3]_net_1 ), 
        .C(\ireg[15]_net_1 ), .Y(\un3_next_sum_m[15] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I149_Y (.A(N621), .B(N625), .Y(
        N702));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I67_Y (.A(N340), .B(N336), .Y(
        N375));
    OR2 next_ireg_3_0_ADD_22x22_fast_I54_Y (.A(N269), .B(I54_un1_Y), 
        .Y(N359));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I378_Y_2 (.A(I118_un1_Y), .B(
        ADD_40x40_fast_I378_Y_0), .C(I194_un1_Y), .Y(
        ADD_40x40_fast_I378_Y_2));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I360_Y (.A(N797), .B(I310_un1_Y), 
        .C(I360_un1_Y), .Y(N1079));
    MX2 \p_adj_RNO[0]  (.A(sr_new[0]), .B(sr_new[0]), .S(sr_new_1_0), 
        .Y(\inf_abs1_5[0] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I384_Y_0 (.A(N691), .B(N684), .C(
        N683), .Y(ADD_40x40_fast_I384_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I182_Y (.A(N658), .B(N655), .C(
        N654), .Y(N735));
    AND3 inf_abs2_a_0_I_52 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[12] ), .Y(N_9_0));
    NOR3A inf_abs2_a_0_I_31 (.A(\DWACT_FINC_E_0[6] ), .B(integral[16]), 
        .C(integral[15]), .Y(N_16));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I232_un1_Y (.A(N717), .B(N710), 
        .Y(I232_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I163_Y (.A(N639), .B(N635), .Y(
        N716));
    NOR3B \ireg_RNIHI7M_0[7]  (.A(\state[3]_net_1 ), .B(
        \ireg[7]_net_1 ), .C(integral[25]), .Y(\ireg_m[7] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I110_Y (.A(N392), .B(N385), .C(
        N384), .Y(N424));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I197_Y (.A(
        ADD_40x40_fast_I197_Y_1), .B(N682), .Y(N756));
    DFN1E1C0 \i_adj[18]  (.D(\inf_abs2_5[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[18]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I91_Y (.A(N511), .B(N508), .Y(
        N641));
    AO1D un1_sumreg_0_0_ADD_40x40_fast_I25_P0N (.A(
        \un1_next_sum_0_iv_1[25] ), .B(\ireg_m[25] ), .C(
        \sumreg[25]_net_1 ), .Y(N547));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I144_Y (.A(N620), .B(N617), .C(
        N616), .Y(N697));
    MX2 \i_adj_RNO[16]  (.A(integral[22]), .B(\inf_abs2_a_0[16] ), .S(
        integral_0_0), .Y(\inf_abs2_5[16] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I71_Y (.A(N538), .B(N541), .Y(
        N621));
    OR3 \ireg_RNIJ2O71[25]  (.A(next_sum_1_sqmuxa_2), .B(
        next_sum_1_sqmuxa_1), .C(\un3_next_sum_m[25] ), .Y(
        \un1_next_sum_0_iv_1[25] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I95_Y (.A(N505), .B(N502), .Y(
        N645));
    OR2 next_ireg_3_0_ADD_22x22_fast_I13_P0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[15]_net_1 ), .Y(N306));
    XA1B \state_RNIGSMMI8[2]  (.A(N1021), .B(ADD_40x40_fast_I457_Y_0), 
        .C(\state[2]_net_1 ), .Y(\next_sum[39] ));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I161_Y (.A(\i_adj[3]_net_1 ), .B(
        \i_adj[1]_net_1 ), .C(N266), .Y(\next_ireg_3[7] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I70_Y (.A(N343), .B(N340), .C(
        N339), .Y(N378));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I75_Y (.A(sum_21), .B(
        \un1_next_sum[21] ), .C(N532), .Y(N625));
    OR3 \ireg_RNIJ45P1[10]  (.A(\un24_next_sum_m[10] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[10] ), .Y(
        \un1_next_sum_iv_2[10] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I168_Y (.A(I168_un1_Y), .B(N640), 
        .Y(N721));
    MX2 \p_adj_RNO[6]  (.A(sr_new[6]), .B(\inf_abs1_a_2[6] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[6] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I379_Y_3 (.A(N756), .B(N771), .C(
        ADD_40x40_fast_I379_Y_2), .Y(ADD_40x40_fast_I379_Y_3));
    OR3 \ireg_RNII03H1[17]  (.A(\un24_next_sum_m[17] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[17] ), .Y(
        \un1_next_sum_iv_2[17] ));
    MX2 \i_adj_RNO[1]  (.A(integral[7]), .B(\inf_abs2_a_0[1] ), .S(
        integral_0_0), .Y(\inf_abs2_5[1] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I75_Y (.A(N344), .B(N348), .Y(
        N383));
    GND GND_i (.Y(GND));
    OR2 next_ireg_3_0_ADD_22x22_fast_I3_P0N (.A(\i_adj[3]_net_1 ), .B(
        \i_adj[5]_net_1 ), .Y(N276));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I143_Y_0 (.A(\i_adj[17]_net_1 ), 
        .B(\i_adj[19]_net_1 ), .C(N314), .Y(ADD_22x22_fast_I143_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I244_un1_Y (.A(N729), .B(N722), 
        .Y(I244_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I348_un1_Y_0 (.A(N790), .B(
        N774), .Y(ADD_40x40_fast_I348_un1_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I244_Y (.A(I244_un1_Y), .B(N721), 
        .Y(N803));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I314_Y (.A(N802), .B(N817), .C(
        N801), .Y(N1085));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I320_Y (.A(N731), .B(I254_un1_Y), 
        .C(I320_un1_Y), .Y(N1103));
    NOR3 \state_RNII1EM[6]  (.A(sum_rdy), .B(\state[6]_net_1 ), .C(
        \state[1]_net_1 ), .Y(\state_RNII1EM[6]_net_1 ));
    MX2 \p_adj_RNO[5]  (.A(sr_new[5]), .B(\inf_abs1_a_2[5] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[5] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I378_Y_3 (.A(N754), .B(N769), .C(
        ADD_40x40_fast_I378_Y_2), .Y(ADD_40x40_fast_I378_Y_3));
    DFN1C0 \state[5]  (.D(\state[4]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[5]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I78_Y (.A(N351), .B(N348), .C(
        N347), .Y(N386));
    NOR2 inf_abs2_a_0_I_21 (.A(integral[12]), .B(integral[13]), .Y(
        \DWACT_FINC_E[3] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I418_Y_0 (.A(sum_0_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I418_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I87_Y (.A(N514), .B(N517), .Y(
        N637));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I29_Y (.A(N306), .B(N309), .Y(
        N334));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I22_P0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[22] ), .C(sum_22), .Y(N538));
    NOR3A inf_abs1_a_2_I_31 (.A(\DWACT_FINC_E[6] ), .B(sr_new[9]), .C(
        sr_new[10]), .Y(N_3));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I27_Y (.A(N309), .B(N312), .Y(
        N332));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I223_Y (.A(N700), .B(N708), .Y(
        N782));
    OR3 \preg_RNIV6PI1[7]  (.A(\un24_next_sum_m[7] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[7] ), .Y(
        \un1_next_sum_iv_2[7] ));
    DFN1E1C0 \ireg[6]  (.D(\next_ireg_3[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[6]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I334_un1_Y (.A(N842), .B(N873), 
        .Y(I334_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I349_un1_Y_0 (.A(N792), .B(
        N776), .Y(ADD_40x40_fast_I349_un1_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I23_G0N (.A(\un1_next_sum[23] )
        , .B(sum_23), .Y(N540));
    DFN1E1C0 \preg[6]  (.D(\p_adj[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[6]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I36_Y (.A(N293), .B(N297), .C(
        N296), .Y(N341));
    NOR2 inf_abs1_a_2_I_6 (.A(sr_new[0]), .B(sr_new[1]), .Y(N_12));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I1_G0N (.A(\i_adj[1]_net_1 ), 
        .B(\i_adj[3]_net_1 ), .Y(N269));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I318_Y (.A(N810), .B(N743), .C(
        N809), .Y(N1097));
    OR2 next_ireg_3_0_ADD_22x22_fast_I114_Y (.A(I114_un1_Y), .B(N390), 
        .Y(N528));
    AO13 un1_sumreg_0_0_ADD_40x40_fast_I64_Y (.A(\sumreg[26]_net_1 ), 
        .B(N546), .C(\un1_next_sum_1_iv[26] ), .Y(N614));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I457_Y_0 (.A(sum_39), .B(
        \un1_next_sum_1_iv[26] ), .Y(ADD_40x40_fast_I457_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I208_un1_Y (.A(N693), .B(N686), 
        .Y(I208_un1_Y));
    XA1B \sumreg_RNO[34]  (.A(N1031), .B(ADD_40x40_fast_I452_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[34] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I81_Y (.A(N354), .B(N350), .Y(
        N389));
    OR2 \ireg_RNILQP41[19]  (.A(\un1_next_sum_iv_0[19] ), .B(
        \un1_next_sum_2[4] ), .Y(\un1_next_sum[19] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I128_Y (.A(N600), .B(N604), .Y(
        N681));
    DFN1E1C0 \sumreg[29]  (.D(\next_sum[29] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[29]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I99_Y (.A(N499), .B(N496), .Y(
        N649));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I169_Y_0 (.A(\i_adj[11]_net_1 ), 
        .B(\i_adj[9]_net_1 ), .Y(ADD_22x22_fast_I169_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I226_Y (.A(N711), .B(N704), .C(
        N703), .Y(N785));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I442_Y_0 (.A(\sumreg[24]_net_1 )
        , .B(\un1_next_sum[24] ), .Y(ADD_40x40_fast_I442_Y_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I212_Y (.A(N608), .B(N612), .C(
        I212_un1_Y), .Y(N771));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I79_Y (.A(N529), .B(N526), .Y(
        N629));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I167_Y (.A(N639), .B(N643), .Y(
        N720));
    NOR3 inf_abs1_a_2_I_10 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2])
        , .Y(\DWACT_FINC_E[0] ));
    DFN1C0 \state_0[3]  (.D(\state[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_0[3]_net_1 ));
    DFN1E1C0 \ireg[21]  (.D(\next_ireg_3[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[21]_net_1 ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I281_Y (.A(N694), .B(N686), .C(
        N784), .Y(N852));
    XNOR2 inf_abs2_a_0_I_32 (.A(integral[17]), .B(N_16), .Y(
        \inf_abs2_a_0[11] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I430_Y_0 (.A(
        \un1_next_sum_iv_1[12] ), .B(\un1_next_sum_iv_2[12] ), .C(
        sum_12), .Y(ADD_40x40_fast_I430_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I217_Y (.A(N694), .B(N702), .Y(
        N776));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I15_P0N (.A(
        \un1_next_sum_iv_1[15] ), .B(\un1_next_sum_iv_2[15] ), .C(
        sum_15), .Y(N517));
    XA1B \sumreg_RNO[27]  (.A(N1049), .B(ADD_40x40_fast_I445_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[27] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I74_Y (.A(N347), .B(N344), .C(
        N343), .Y(N382));
    DFN1E1C0 \sumreg[19]  (.D(\next_sum[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_19));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I422_Y_0 (.A(
        \un1_next_sum_2[4] ), .B(\un1_next_sum_iv_0[4] ), .C(sum_4), 
        .Y(ADD_40x40_fast_I422_Y_0));
    DFN1E1C0 \sumreg[8]  (.D(\next_sum[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_8));
    NOR2A \state_RNIBU9J_0[3]  (.A(\state[3]_net_1 ), .B(integral[25]), 
        .Y(next_sum_1_sqmuxa));
    DFN1E1C0 \sumreg[28]  (.D(\next_sum[28] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[28]_net_1 ));
    XA1B \sumreg_RNO[0]  (.A(N_228), .B(ADD_40x40_fast_I418_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[0] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I430_Y (.A(
        ADD_40x40_fast_I430_Y_0), .B(N1094), .Y(\un1_sumreg[12] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I256_un1_Y (.A(N741), .B(N734), 
        .Y(I256_un1_Y));
    NOR3B \ireg_RNIHI7M[7]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[7]_net_1 ), .Y(\un3_next_sum_m[7] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I451_Y_0 (.A(
        \sumreg[33]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I451_Y_0));
    AO1 un1_sumreg_0_0_ADD_m8_i_1 (.A(ADD_m8_i_a4_0_1), .B(N_232), .C(
        \un1_next_sum_2[4] ), .Y(ADD_m8_i_1));
    AO1 \ireg_RNIHNU91[14]  (.A(\ireg[14]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[14] ), .Y(
        \un1_next_sum_iv_1[14] ));
    OR2 \ireg_RNIHNQ41[24]  (.A(\un1_next_sum_iv_0[24] ), .B(
        \un1_next_sum_2[4] ), .Y(\un1_next_sum[24] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I143_Y (.A(N615), .B(N619), .Y(
        N696));
    NOR3A \state_RNIPCJR[4]  (.A(integral_0_0), .B(\state[5]_net_1 ), 
        .C(\state[4]_net_1 ), .Y(N_232));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_1_0 (.A(
        ADD_22x22_fast_I142_Y_0_a3_0), .B(N330), .Y(
        ADD_22x22_fast_I142_Y_0_a3_1));
    DFN1C0 \state_2[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_2[2]_net_1 ));
    DFN1E1C0 \sumreg[18]  (.D(\next_sum[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_18));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I380_Y_1 (.A(I122_un1_Y), .B(
        N594), .C(N683), .Y(ADD_40x40_fast_I380_Y_1));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I61_Y (.A(\sumreg[27]_net_1 ), 
        .B(\sumreg[28]_net_1 ), .C(\un1_next_sum_1_iv[26] ), .Y(N611));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I6_G0N (.A(\i_adj[6]_net_1 ), 
        .B(\i_adj[8]_net_1 ), .Y(N284));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I162_Y (.A(\i_adj[4]_net_1 ), .B(
        \i_adj[2]_net_1 ), .C(N359), .Y(\next_ireg_3[8] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I243_Y (.A(N728), .B(N720), .Y(
        N802));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I127_Y (.A(N599), .B(N603), .Y(
        N680));
    DFN1E1C0 \p_adj[3]  (.D(\inf_abs1_5[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[3]_net_1 ));
    DFN1E1C0 \ireg[10]  (.D(\next_ireg_3[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[10]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I49_Y (.A(N276), .B(N279), .Y(
        N354));
    OA1A un1_sumreg_0_0_ADD_40x40_fast_I65_Y (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[26]_net_1 ), .C(N547), .Y(
        N615));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I47_Y (.A(N279), .B(N282), .Y(
        N352));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I101_Y (.A(N496), .B(N493), .Y(
        N651));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I12_P0N (.A(
        \un1_next_sum_iv_1[12] ), .B(\un1_next_sum_iv_2[12] ), .C(
        sum_12), .Y(N508));
    NOR2B \ireg_RNI18LJ[25]  (.A(\ireg[25]_net_1 ), .B(
        next_sum_0_sqmuxa), .Y(\ireg_m[25] ));
    AND3 inf_abs2_a_0_I_22 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_19));
    DFN1E1C0 \sumreg[1]  (.D(\next_sum[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_1_d0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I131_un1_Y_0 (.A(N389), .B(N381)
        , .Y(ADD_22x22_fast_I131_un1_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I449_Y_0 (.A(
        \sumreg[31]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I449_Y_0));
    XA1B \sumreg_RNO[20]  (.A(N1070), .B(ADD_40x40_fast_I438_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[20] ));
    DFN1E1C0 \sumreg_0[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(sum_0_0));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I47_Y (.A(\sumreg[35]_net_1 ), 
        .B(\sumreg[34]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N597)
        );
    XNOR2 inf_abs1_a_2_I_32 (.A(sr_new[11]), .B(N_3), .Y(
        \inf_abs1_a_2[11] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I187_Y_0 (.A(sum_1_d0), .B(
        sum_2_d0), .C(\un1_next_sum[0] ), .Y(ADD_40x40_fast_I187_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I148_Y (.A(N624), .B(N621), .C(
        N620), .Y(N701));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I165_Y (.A(
        ADD_22x22_fast_I165_Y_0), .B(N531), .Y(\next_ireg_3[11] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I13_G0N (.A(
        \un1_next_sum_iv_1[13] ), .B(\un1_next_sum_iv_2[13] ), .C(
        sum_13), .Y(N510));
    XA1B \sumreg_RNO[21]  (.A(N1067), .B(ADD_40x40_fast_I439_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[21] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_3_0 (.A(N338), .B(
        N334), .Y(ADD_22x22_fast_I142_Y_0_a3_3_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I131_Y (.A(N607), .B(N603), .Y(
        N684));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I303_Y (.A(N806), .B(N790), .Y(
        N874));
    XNOR2 inf_abs1_a_2_I_20 (.A(sr_new[7]), .B(N_7_0), .Y(
        \inf_abs1_a_2[7] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I438_Y_0 (.A(sum_20), .B(
        \un1_next_sum[20] ), .Y(ADD_40x40_fast_I438_Y_0));
    DFN1E1C0 \sumreg[25]  (.D(\next_sum[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[25]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I246_Y (.A(N731), .B(N724), .C(
        N723), .Y(N805));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I151_Y (.A(N623), .B(N627), .Y(
        N704));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I176_Y (.A(N652), .B(N649), .C(
        N648), .Y(N729));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I347_Y (.A(
        ADD_40x40_fast_I347_un1_Y_0), .B(N1088), .C(
        ADD_40x40_fast_I347_Y_0), .Y(N1040));
    NOR3B \preg_RNI2IN01[14]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), 
        .C(\preg[14]_net_1 ), .Y(\un24_next_sum_m[14] ));
    DFN1E1C0 \ireg[23]  (.D(\next_ireg_3[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[23]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I106_un1_Y (.A(N381), .B(N388), 
        .Y(I106_un1_Y));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I429_Y_0 (.A(sum_11), .B(
        \un1_next_sum[11] ), .Y(ADD_40x40_fast_I429_Y_0));
    OR2 un1_sumreg_0_0_ADD_m8_i (.A(ADD_m8_i_1), .B(ADD_m8_i_a4_3), .Y(
        N743));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I9_G0N (.A(\un1_next_sum[9] ), 
        .B(sum_9), .Y(N498_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I447_Y_0 (.A(
        \sumreg[29]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I447_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I353_Y (.A(
        ADD_40x40_fast_I353_un1_Y_0), .B(N1106), .C(
        ADD_40x40_fast_I353_Y_0), .Y(N1058));
    NOR3B \preg_RNIVEN01[11]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), 
        .C(\preg[11]_net_1 ), .Y(\un24_next_sum_m[11] ));
    NOR3B \ireg_RNIQMMG_0[10]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[10]_net_1 ), .C(integral_1_0), .Y(\ireg_m[10] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I379_Y_4 (.A(N840), .B(N871), .C(
        ADD_40x40_fast_I379_Y_3), .Y(ADD_40x40_fast_I379_Y_4));
    AO1 \preg_RNINDR41[8]  (.A(\preg[8]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[8] ), .Y(
        \un1_next_sum_iv_1[8] ));
    AND3 inf_abs2_a_0_I_60 (.A(integral_i[24]), .B(integral_i[25]), .C(
        integral_i[25]), .Y(\DWACT_FINC_E[15] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I170_Y (.A(N646), .B(N643), .C(
        N642), .Y(N723));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I166_un1_Y (.A(N642), .B(N639), 
        .Y(I166_un1_Y));
    OR3 \state_RNITOC71_0[4]  (.A(next_sum_1_sqmuxa_2), .B(
        next_sum_1_sqmuxa_1), .C(next_sum_1_sqmuxa), .Y(
        \un1_next_sum_1_iv[26] ));
    NOR3B \ireg_RNIHAK8[16]  (.A(integral_1_0), .B(\state[3]_net_1 ), 
        .C(\ireg[16]_net_1 ), .Y(\un3_next_sum_m[16] ));
    DFN1E1C0 \sumreg[15]  (.D(\next_sum[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_15));
    DFN1E1C0 \ireg[5]  (.D(\i_adj[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[5]_net_1 ));
    DFN1E1C0 \ireg[25]  (.D(\next_ireg_3[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[25]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0 (.A(
        ADD_22x22_fast_I142_Y_0_a3_1), .B(N_11), .C(
        ADD_22x22_fast_I142_Y_0_1), .Y(N492));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I353_Y_0 (.A(N799), .B(N784), .C(
        N783), .Y(ADD_40x40_fast_I353_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I5_G0N (.A(\un1_next_sum[5] ), 
        .B(sum_5), .Y(N486));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I427_Y_0 (.A(sum_9), .B(
        \un1_next_sum[9] ), .Y(ADD_40x40_fast_I427_Y_0));
    DFN1E1C0 \p_adj[9]  (.D(\inf_abs1_5[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[9]_net_1 ));
    XNOR2 inf_abs1_a_2_I_17 (.A(sr_new[6]), .B(N_8_0), .Y(
        \inf_abs1_a_2[6] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I163_Y (.A(
        ADD_22x22_fast_I163_Y_0), .B(N396), .Y(\next_ireg_3[9] ));
    OR2 \state_RNITOC71[3]  (.A(\un1_next_sum_2[4] ), .B(
        next_sum_0_sqmuxa), .Y(\un1_next_sum[0] ));
    MX2 \i_adj_RNO[14]  (.A(integral[20]), .B(\inf_abs2_a_0[14] ), .S(
        integral_0_0), .Y(\inf_abs2_5[14] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I69_Y (.A(N544), .B(N541), .Y(
        N619));
    XA1B \sumreg_RNO[14]  (.A(N1088), .B(ADD_40x40_fast_I432_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[14] ));
    XA1B \sumreg_RNO[35]  (.A(N1029), .B(ADD_40x40_fast_I453_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[35] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I349_Y (.A(
        ADD_40x40_fast_I349_un1_Y_0), .B(N1094), .C(
        ADD_40x40_fast_I349_Y_0), .Y(N1046));
    NOR3B \ireg_RNIF8K8[14]  (.A(integral_1_0), .B(\state[3]_net_1 ), 
        .C(\ireg[14]_net_1 ), .Y(\un3_next_sum_m[14] ));
    DFN1C0 \state[4]  (.D(\state_0[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[4]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I147_Y (.A(N623), .B(N619), .Y(
        N700));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I8_G0N (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[8]_net_1 ), .Y(N290));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_0 (.A(\i_adj[18]_net_1 )
        , .B(\i_adj[20]_net_1 ), .C(N_14_1), .Y(
        ADD_22x22_fast_I142_Y_0_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I9_P0N (.A(\i_adj[9]_net_1 ), .B(
        \i_adj[11]_net_1 ), .Y(N294));
    DFN1E1C0 \sumreg[26]  (.D(\next_sum[26] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[26]_net_1 ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I441_Y_0 (.A(sum_23), .B(
        \un1_next_sum[23] ), .Y(ADD_40x40_fast_I441_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I179_Y (.A(N655), .B(N651), .Y(
        N732));
    XA1B \sumreg_RNO[7]  (.A(N817), .B(ADD_40x40_fast_I425_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[7] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I11_P0N (.A(\un1_next_sum[11] ), 
        .B(sum_11), .Y(N505));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I267_Y (.A(N754), .B(N770), .Y(
        N838));
    AO1 next_ireg_3_0_ADD_22x22_fast_I128_Y_0 (.A(N382), .B(N375), .C(
        N374), .Y(ADD_22x22_fast_I128_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I90_Y (.A(N507_0), .B(N511), .C(
        N510), .Y(N640));
    DFN1E1C0 \ireg[17]  (.D(\next_ireg_3[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[17]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I316_Y (.A(N806), .B(N821), .C(
        N805), .Y(N1091));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I305_Y (.A(N808), .B(N792), .Y(
        N876));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I381_Y (.A(
        ADD_40x40_fast_I381_Y_2), .B(I381_un1_Y), .C(I336_un1_Y), .Y(
        N1027));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I219_Y (.A(N696), .B(N704), .Y(
        N778));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I102_Y (.A(N489), .B(N493), .C(
        N492_0), .Y(N652));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I257_Y_0 (.A(\un1_next_sum[0] ), 
        .B(sum_1_d0), .C(N472), .Y(ADD_40x40_fast_I257_Y_0));
    NOR3C un1_sumreg_0_0_ADD_m8_i_a4_0_1 (.A(sum_1_d0), .B(sum_0_d0), 
        .C(sum_2_d0), .Y(ADD_m8_i_a4_0_1));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I70_Y (.A(N537), .B(N541), .C(
        N540), .Y(N620));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I21_G0N (.A(\un1_next_sum[21] )
        , .B(sum_21), .Y(N534));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I195_Y (.A(N595), .B(N591), .C(
        N680), .Y(N754));
    XA1 \ireg_RNITQNG[22]  (.A(integral_1_0), .B(\ireg[22]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[22] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I421_Y_0 (.A(sum_3), .B(N743), 
        .Y(ADD_40x40_fast_I421_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I174_Y (.A(N650), .B(N647), .C(
        N646), .Y(N727));
    NOR2A \state_RNIRVM7_0[4]  (.A(\state[4]_net_1 ), .B(derivative_0), 
        .Y(next_sum_1_sqmuxa_1));
    DFN1E1C0 \sumreg[16]  (.D(\next_sum[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_16));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I16_G0N (.A(\i_adj[16]_net_1 ), 
        .B(\i_adj[18]_net_1 ), .Y(N314));
    XNOR2 inf_abs2_a_0_I_14 (.A(integral[11]), .B(N_22), .Y(
        \inf_abs2_a_0[5] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I355_Y (.A(I355_un1_Y), .B(N871), 
        .Y(N1064));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I132_Y (.A(N608), .B(N604), .Y(
        N685));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I2_G0N (.A(\i_adj[2]_net_1 ), 
        .B(\i_adj[4]_net_1 ), .Y(N272));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I152_Y (.A(N628), .B(N625), .C(
        N624), .Y(N705));
    MX2 \p_adj_RNO[8]  (.A(sr_new[8]), .B(\inf_abs1_a_2[8] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[8] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I3_P0N (.A(sum_3), .B(
        \un1_next_sum[0] ), .Y(N481));
    AO1 next_ireg_3_0_ADD_22x22_fast_I76_Y (.A(N349), .B(N346), .C(
        N345), .Y(N384));
    DFN1E1C0 \sumreg[21]  (.D(\next_sum[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(sum_21));
    MX2 \p_adj_RNO[7]  (.A(sr_new[7]), .B(\inf_abs1_a_2[7] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[7] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I84_Y (.A(N516), .B(N520), .C(
        N519), .Y(N634));
    AO1 next_ireg_3_0_ADD_22x22_fast_I42_Y (.A(N284), .B(N288), .C(
        N287), .Y(N347));
    NOR3B \ireg_RNITPMG_0[13]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[13]_net_1 ), .C(integral_1_0), .Y(\ireg_m[13] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I222_Y (.A(N707), .B(N700), .C(
        N699), .Y(N781));
    XA1B \sumreg_RNO[36]  (.A(N1027), .B(ADD_40x40_fast_I454_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[36] ));
    NOR2B \preg_RNIJJAM[15]  (.A(\preg[15]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[15] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I31_Y (.A(N303), .B(N306), .Y(
        N336));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I310_un1_Y (.A(N731), .B(
        I254_un1_Y), .C(N798), .Y(I310_un1_Y));
    AO1 next_ireg_3_0_ADD_22x22_fast_I129_Y (.A(
        ADD_22x22_fast_I129_un1_Y_0), .B(N531), .C(
        ADD_22x22_fast_I129_Y_0), .Y(N507));
    NOR3B \ireg_RNIIJ7M_0[8]  (.A(\state[3]_net_1 ), .B(
        \ireg[8]_net_1 ), .C(integral[25]), .Y(\ireg_m[8] ));
    AO1 \ireg_RNIBHU91[11]  (.A(\ireg[11]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[11] ), .Y(
        \un1_next_sum_iv_1[11] ));
    DFN1E1C0 \p_adj[1]  (.D(\inf_abs1_5[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[1]_net_1 ));
    NOR3A inf_abs1_a_2_I_27 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .C(
        sr_new[9]), .Y(N_4));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I186_Y (.A(N662), .B(N659), .C(
        N658), .Y(N739));
    NOR2 inf_abs2_a_0_I_15 (.A(integral[9]), .B(integral[10]), .Y(
        \DWACT_FINC_E[1] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I434_Y_0 (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(ADD_40x40_fast_I434_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I227_Y (.A(N704), .B(N712), .Y(
        N786));
    DFN1E1C0 \p_adj[7]  (.D(\inf_abs1_5[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[7]_net_1 ));
    DFN1E1C0 \sumreg[11]  (.D(\next_sum[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_11));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I433_Y_0 (.A(
        \un1_next_sum_iv_1[15] ), .B(\un1_next_sum_iv_2[15] ), .C(
        sum_15), .Y(ADD_40x40_fast_I433_Y_0));
    XA1B \sumreg_RNO[33]  (.A(N1033), .B(ADD_40x40_fast_I451_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[33] ));
    DFN1E1C0 \ireg[19]  (.D(\next_ireg_3[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[19]_net_1 ));
    NOR2B \state_RNIRVM7[4]  (.A(\state[4]_net_1 ), .B(derivative_0), 
        .Y(next_sum_0_sqmuxa_1));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I320_un1_Y (.A(N814), .B(N666), 
        .Y(I320_un1_Y));
    MX2 \i_adj_RNO[10]  (.A(integral[16]), .B(\inf_abs2_a_0[10] ), .S(
        integral_0_0), .Y(\inf_abs2_5[10] ));
    XNOR2 inf_abs2_a_0_I_40 (.A(integral[20]), .B(N_13), .Y(
        \inf_abs2_a_0[14] ));
    AND3 inf_abs2_a_0_I_54 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E[9] ), .C(\DWACT_FINC_E[12] ), .Y(
        \DWACT_FINC_E[13] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I180_Y (.A(N656), .B(N653), .C(
        N652), .Y(N733));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I167_Y (.A(\i_adj[9]_net_1 ), .B(
        \i_adj[7]_net_1 ), .C(N525), .Y(\next_ireg_3[13] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I57_Y (.A(\sumreg[30]_net_1 ), 
        .B(\sumreg[29]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N607)
        );
    DFN1C0 \state[1]  (.D(\state_RNIAMDD[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[1]_net_1 ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I382_Y (.A(
        ADD_40x40_fast_I382_Y_1), .B(I382_un1_Y), .C(I338_un1_Y), .Y(
        N1029));
    MX2 \p_adj_RNO[10]  (.A(sr_new[10]), .B(\inf_abs1_a_2[10] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[10] ));
    DFN1E1C0 \ireg[22]  (.D(\next_ireg_3[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[22]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I20_P0N (.A(\un1_next_sum[20] ), 
        .B(sum_20), .Y(N532));
    AX1D next_ireg_3_0_ADD_22x22_fast_I169_Y (.A(N424), .B(I133_un1_Y), 
        .C(ADD_22x22_fast_I169_Y_0), .Y(\next_ireg_3[15] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I114_un1_Y (.A(N391), .B(N359), 
        .Y(I114_un1_Y));
    NOR3B inf_abs2_a_0_I_16 (.A(\DWACT_FINC_E[1] ), .B(
        \DWACT_FINC_E_0[0] ), .C(integral[11]), .Y(N_21));
    NOR3B \preg_RNIFFAM[11]  (.A(\state[5]_net_1 ), .B(
        \preg[11]_net_1 ), .C(sr_new[12]), .Y(\preg_m[11] ));
    NOR3B inf_abs2_a_0_I_55 (.A(\DWACT_FINC_E[13] ), .B(
        \DWACT_FINC_E[28] ), .C(integral[24]), .Y(N_8));
    DFN1E1C0 \preg[13]  (.D(\p_adj[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[13]_net_1 ));
    DFN1E1C0 \i_adj[6]  (.D(\inf_abs2_5[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[6]_net_1 ));
    DFN1E1C0 \i_adj[4]  (.D(\inf_abs2_5[4] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[4]_net_1 ));
    NOR2B \state_RNINQBC[5]  (.A(\state[5]_net_1 ), .B(sr_new[12]), .Y(
        next_sum_0_sqmuxa_2));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I63_Y (.A(N332), .B(N336), .Y(
        N371));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I230_Y (.A(N715), .B(N708), .C(
        N707), .Y(N789));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I81_Y (.A(N526), .B(N523), .Y(
        N631));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I379_Y_2 (.A(N596), .B(
        ADD_40x40_fast_I379_Y_0), .C(N681), .Y(ADD_40x40_fast_I379_Y_2)
        );
    MX2 \i_adj_RNO[18]  (.A(integral[24]), .B(\inf_abs2_a_0[18] ), .S(
        integral_0_0), .Y(\inf_abs2_5[18] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I250_Y (.A(N735), .B(N728), .C(
        N727), .Y(N809));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I456_Y_0 (.A(
        \sumreg[38]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I456_Y_0));
    NOR2A inf_abs1_a_2_I_11 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .Y(
        N_10));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I348_Y (.A(
        ADD_40x40_fast_I348_un1_Y_0), .B(N1091), .C(
        ADD_40x40_fast_I348_Y_0), .Y(N1043));
    OR2 \preg_RNIDJHS[6]  (.A(next_sum_0_sqmuxa_1), .B(
        \un24_next_sum_m[6] ), .Y(\un1_next_sum_iv_0[6] ));
    NOR3B \preg_RNI6MN01[18]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), 
        .C(\preg[18]_net_1 ), .Y(\un24_next_sum_m[18] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I381_Y_1 (.A(N596), .B(N600), .C(
        N685), .Y(ADD_40x40_fast_I381_Y_1));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I92_Y (.A(N504_0), .B(N508), .C(
        N507_0), .Y(N642));
    DFN1E1C0 \i_adj[9]  (.D(\inf_abs2_5[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[9]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I85_Y (.A(N517), .B(N520), .Y(
        N635));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I11_G0N (.A(\un1_next_sum[11] )
        , .B(sum_11), .Y(N504_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I201_Y (.A(
        ADD_40x40_fast_I201_Y_0), .B(N686), .Y(N760));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I72_Y (.A(N534), .B(N538), .C(
        N537), .Y(N622));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I0_S (.A(\i_adj[0]_net_1 ), .B(
        \i_adj[2]_net_1 ), .Y(\next_ireg_3[6] ));
    NOR3B \preg_RNILMQK[9]  (.A(sr_new_0_0), .B(\state[5]_net_1 ), .C(
        \preg[9]_net_1 ), .Y(\un24_next_sum_m[9] ));
    DFN1E1C0 \i_adj[3]  (.D(\inf_abs2_5[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[3]_net_1 ));
    XA1B \sumreg_RNO[15]  (.A(N1085), .B(ADD_40x40_fast_I433_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[15] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I242_Y (.A(N727), .B(N720), .C(
        N719), .Y(N801));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y_1 (.A(N371), .B(N378), .C(
        ADD_22x22_fast_I126_Y_0), .Y(ADD_22x22_fast_I126_Y_1));
    OR2 next_ireg_3_0_ADD_22x22_fast_I14_P0N (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .Y(N309));
    OA1 next_ireg_3_0_ADD_22x22_fast_I51_Y (.A(\i_adj[4]_net_1 ), .B(
        \i_adj[2]_net_1 ), .C(N276), .Y(N356));
    AX1D next_ireg_3_0_ADD_22x22_fast_I178_Y (.A(I122_un1_Y_0), .B(
        ADD_22x22_fast_I143_Y_3), .C(ADD_22x22_fast_I178_Y_0), .Y(
        \next_ireg_3[24] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I231_Y (.A(N716), .B(N708), .Y(
        N790));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I184_Y (.A(N660), .B(N657), .C(
        N656), .Y(N737));
    XNOR2 inf_abs2_a_0_I_56 (.A(integral[25]), .B(N_8), .Y(
        \inf_abs2_a_0[19] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I87_Y (.A(I54_un1_Y), .B(N357), 
        .Y(N396));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I251_Y (.A(N736), .B(N728), .Y(
        N810));
    DFN1E1C0 \sumreg[34]  (.D(\next_sum[34] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[34]_net_1 ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I340_un1_Y (.A(N795), .B(
        I308_un1_Y), .C(N848), .Y(I340_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I247_Y (.A(N724), .B(N732), .Y(
        N806));
    DFN1C0 \state_0[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_0[2]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I60_Y (.A(\sumreg[27]_net_1 ), 
        .B(\sumreg[28]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N610)
        );
    OR3 \ireg_RNIPA5P1[13]  (.A(\un24_next_sum_m[13] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[13] ), .Y(
        \un1_next_sum_iv_2[13] ));
    AO1 \preg_RNIPFR41[9]  (.A(\preg[9]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[9] ), .Y(
        \un1_next_sum_iv_1[9] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I385_un1_Y (.A(N884), .B(
        \un1_next_sum[0] ), .C(N852), .Y(I385_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I173_Y (.A(N645), .B(N649), .Y(
        N726));
    DFN1E1C0 \ireg[7]  (.D(\next_ireg_3[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[7]_net_1 ));
    XA1B \sumreg_RNO[28]  (.A(N1046), .B(ADD_40x40_fast_I446_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[28] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I380_un1_Y (.A(N821), .B(N874), 
        .C(N842), .Y(I380_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I238_Y (.A(N723), .B(N716), .C(
        N715), .Y(N797));
    XA1B \sumreg_RNO[3]  (.A(\un1_next_sum[0] ), .B(
        ADD_40x40_fast_I421_Y_0), .C(\state[2]_net_1 ), .Y(
        \next_sum[3] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I269_Y (.A(N756), .B(N772), .Y(
        N840));
    DFN1E1C0 \preg[7]  (.D(\p_adj[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[7]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I44_Y (.A(\sumreg[35]_net_1 ), 
        .B(\sumreg[36]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N594)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I258_Y (.A(N736), .B(N743), .C(
        N735), .Y(N817));
    NOR3B \preg_RNI5LN01[17]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), 
        .C(\preg[17]_net_1 ), .Y(\un24_next_sum_m[17] ));
    OR3 next_ireg_3_0_ADD_22x22_fast_I131_Y (.A(I131_un1_Y), .B(
        ADD_22x22_fast_I131_Y_0), .C(I106_un1_Y), .Y(N513));
    DFN1E1C0 \ireg[16]  (.D(\next_ireg_3[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[16]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I273_Y (.A(N760), .B(N776), .Y(
        N844));
    OR2 \state_RNIIQ2K[5]  (.A(next_sum_0_sqmuxa_1), .B(
        next_sum_0_sqmuxa_2), .Y(\un1_next_sum_2[4] ));
    XA1B \sumreg_RNO[32]  (.A(N1035), .B(ADD_40x40_fast_I450_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[32] ));
    DFN1E1C0 \preg[10]  (.D(\p_adj[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[10]_net_1 ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I163_Y_0 (.A(\i_adj[5]_net_1 ), 
        .B(\i_adj[3]_net_1 ), .Y(ADD_22x22_fast_I163_Y_0));
    AO1 \ireg_RNIPVU91[18]  (.A(\ireg[18]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[18] ), .Y(
        \un1_next_sum_iv_1[18] ));
    DFN1E1C0 \preg[18]  (.D(\p_adj[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[18]_net_1 ));
    NOR3 inf_abs2_a_0_I_18 (.A(integral[10]), .B(integral[9]), .C(
        integral[11]), .Y(\DWACT_FINC_E[2] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I6_P0N (.A(\un1_next_sum[6] ), 
        .B(sum_6), .Y(N490));
    XA1B \sumreg_RNO[8]  (.A(N1106), .B(ADD_40x40_fast_I426_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[8] ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I23_Y (.A(\i_adj[18]_net_1 ), .B(
        \i_adj[16]_net_1 ), .C(N_9), .Y(N328));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I178_Y (.A(N654), .B(N651), .C(
        N650), .Y(N731));
    NOR2B inf_abs2_a_0_I_34 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .Y(N_15));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I98_Y (.A(N495), .B(N499), .C(
        N498_0), .Y(N648));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I7_P0N (.A(\un1_next_sum[7] ), 
        .B(sum_7), .Y(N493));
    NOR2 inf_abs2_a_0_I_47 (.A(integral[21]), .B(integral[22]), .Y(
        \DWACT_FINC_E[11] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I89_Y (.A(N514), .B(N511), .Y(
        N639));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I10_P0N (.A(
        \un1_next_sum_iv_1[10] ), .B(\un1_next_sum_iv_2[10] ), .C(
        sum_10), .Y(N502));
    NOR2 inf_abs1_a_2_I_21 (.A(sr_new[6]), .B(sr_new[7]), .Y(
        \DWACT_FINC_E_0[3] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I5_G0N (.A(\i_adj[5]_net_1 ), 
        .B(\i_adj[7]_net_1 ), .Y(N281));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I176_Y (.A(\i_adj[16]_net_1 ), 
        .B(\i_adj[18]_net_1 ), .C(N498), .Y(\next_ireg_3[22] ));
    NOR3 inf_abs2_a_0_I_8 (.A(integral[7]), .B(integral[6]), .C(
        integral[8]), .Y(N_24));
    XA1B \sumreg_RNO[16]  (.A(N1082), .B(ADD_40x40_fast_I434_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[16] ));
    NOR3B inf_abs2_a_0_I_19 (.A(\DWACT_FINC_E[2] ), .B(
        \DWACT_FINC_E_0[0] ), .C(integral[12]), .Y(N_20));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I78_Y (.A(N525_0), .B(N529), .C(
        N528_0), .Y(N628));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I132_un1_Y (.A(N423), .B(N359), 
        .Y(I132_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I0_CO1 (.A(\i_adj[0]_net_1 ), 
        .B(\i_adj[2]_net_1 ), .Y(N266));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I229_Y (.A(N706), .B(N714), .Y(
        N788));
    XA1B \sumreg_RNO[13]  (.A(N1091), .B(ADD_40x40_fast_I431_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[13] ));
    XA1 \ireg_RNI30NG[19]  (.A(integral_1_0), .B(\ireg[19]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[19] ));
    XNOR2 inf_abs2_a_0_I_7 (.A(integral[8]), .B(N_25), .Y(
        \inf_abs2_a_0[2] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I133_un1_Y (.A(N425), .B(N266), 
        .Y(I133_un1_Y));
    XNOR2 inf_abs2_a_0_I_35 (.A(integral[18]), .B(N_15), .Y(
        \inf_abs2_a_0[12] ));
    OR3 \ireg_RNIL65P1[11]  (.A(\un24_next_sum_m[11] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[11] ), .Y(
        \un1_next_sum_iv_2[11] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I1_P0N (.A(\i_adj[1]_net_1 ), .B(
        \i_adj[3]_net_1 ), .Y(N270));
    XOR2 inf_abs2_a_0_I_5 (.A(integral[6]), .B(integral[7]), .Y(
        \inf_abs2_a_0[1] ));
    AND3 inf_abs2_a_0_I_61 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[15] ), .Y(N_6));
    AND3 inf_abs2_a_0_I_58 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[14] ), .Y(N_7));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I111_Y (.A(\un1_next_sum[0] ), 
        .B(sum_2_d0), .C(N481), .Y(N661));
    XA1B \sumreg_RNO[19]  (.A(N1073), .B(ADD_40x40_fast_I437_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[19] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I68_Y (.A(N341), .B(N338), .C(
        N337), .Y(N376));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I16_G0N (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(N519));
    XNOR2 inf_abs1_a_2_I_12 (.A(sr_new[4]), .B(N_10), .Y(
        \inf_abs1_a_2[4] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I41_Y (.A(\sumreg[38]_net_1 ), 
        .B(\sumreg[37]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N591)
        );
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I446_Y_0 (.A(
        \sumreg[28]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I446_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I109_Y (.A(N391), .B(N383), .Y(
        N423));
    NOR3B \ireg_RNI0L7B[6]  (.A(integral_1_0), .B(\state[3]_net_1 ), 
        .C(\ireg[6]_net_1 ), .Y(\un3_next_sum_m[6] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I93_Y (.A(N508), .B(N505), .Y(
        N643));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I212_un1_Y (.A(N697), .B(N690), 
        .Y(I212_un1_Y));
    DFN1E1C0 \p_adj[12]  (.D(\inf_abs1_5[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[12]_net_1 ));
    DFN1E1C0 \p_adj[2]  (.D(\inf_abs1_5[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[2]_net_1 ));
    MX2 \i_adj_RNO[9]  (.A(integral[15]), .B(\inf_abs2_a_0[9] ), .S(
        integral_0_0), .Y(\inf_abs2_5[9] ));
    DFN1E1C0 \ireg[18]  (.D(\next_ireg_3[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[18]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_1 (.A(N328), .B(N331), .C(
        ADD_22x22_fast_I143_Y_0), .Y(ADD_22x22_fast_I143_Y_1));
    NOR3A inf_abs2_a_0_I_13 (.A(\DWACT_FINC_E_0[0] ), .B(integral[9]), 
        .C(integral[10]), .Y(N_22));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I313_Y (.A(N734), .B(
        ADD_40x40_fast_I257_Y_1), .C(N800), .Y(N884));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I73_Y (.A(sum_21), .B(
        \un1_next_sum[21] ), .C(N538), .Y(N623));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_3 (.A(
        ADD_22x22_fast_I143_un1_Y_0), .B(N423), .C(
        ADD_22x22_fast_I143_Y_2), .Y(ADD_22x22_fast_I143_Y_3));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I45_Y (.A(\sumreg[36]_net_1 ), 
        .B(\sumreg[35]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N595)
        );
    DFN1E1C0 \ireg[9]  (.D(\next_ireg_3[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[9]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I382_Y_0 (.A(I194_un1_Y), .B(
        N687), .Y(ADD_40x40_fast_I382_Y_0));
    DFN1E1C0 \preg[14]  (.D(\p_adj[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[14]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I96_Y (.A(N498_0), .B(N502), .C(
        N501), .Y(N646));
    XNOR2 inf_abs2_a_0_I_59 (.A(integral[25]), .B(N_7), .Y(
        \inf_abs2_a_0[20] ));
    AND3 inf_abs2_a_0_I_24 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E_0[4] ));
    OR2 \state_RNIB7MF1[4]  (.A(N_232), .B(\un1_next_sum_2[4] ), .Y(
        N_228));
    DFN1E1C0 \preg[9]  (.D(\p_adj[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[9]_net_1 ));
    OR2 \ireg_RNI3BPI1[9]  (.A(\un3_next_sum_m[9] ), .B(
        \un1_next_sum_iv_0[9] ), .Y(\un1_next_sum_iv_2[9] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I426_Y_0 (.A(
        \un1_next_sum_iv_1[8] ), .B(\un1_next_sum_iv_2[8] ), .C(sum_8), 
        .Y(ADD_40x40_fast_I426_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I379_Y (.A(
        ADD_40x40_fast_I379_un1_Y_0), .B(N819), .C(
        ADD_40x40_fast_I379_Y_4), .Y(N1023));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I76_Y (.A(N528_0), .B(N532), .C(
        N531_0), .Y(N626));
    DFN1P0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .PRE(n_rst_c), 
        .Q(sum_rdy));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I205_Y (.A(N690), .B(N682), .Y(
        N764));
    NOR2B inf_abs1_a_2_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_2));
    NOR3B inf_abs2_a_0_I_36 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .C(integral[18]), .Y(N_14));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I8_G0N (.A(
        \un1_next_sum_iv_1[8] ), .B(\un1_next_sum_iv_2[8] ), .C(sum_8), 
        .Y(N495));
    XA1B \sumreg_RNO[6]  (.A(N819), .B(ADD_40x40_fast_I424_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[6] ));
    NOR3B \preg_RNI0GN01[12]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), 
        .C(\preg[12]_net_1 ), .Y(\un24_next_sum_m[12] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I71_Y (.A(N344), .B(N340), .Y(
        N379));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I145_Y (.A(N617), .B(N621), .Y(
        N698));
    AO1A \state_RNO[0]  (.A(sum_enable), .B(sum_rdy), .C(
        \state[5]_net_1 ), .Y(\state_ns[0] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I62_Y (.A(\sumreg[26]_net_1 ), 
        .B(\sumreg[27]_net_1 ), .C(\un1_next_sum_1_iv[26] ), .Y(N612));
    OR2 \ireg_RNI01D71[5]  (.A(\un1_next_sum_iv_0[5] ), .B(
        \un1_next_sum_2[4] ), .Y(\un1_next_sum[5] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I380_Y (.A(I380_un1_Y), .B(
        ADD_40x40_fast_I380_Y_2), .C(I334_un1_Y), .Y(N1025));
    NOR3B \ireg_RNIIJ7M[8]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[8]_net_1 ), .Y(\un3_next_sum_m[8] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I235_Y (.A(N712), .B(N720), .Y(
        N794));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I191_Y (.A(I116_un1_Y), .B(N664), 
        .Y(N745));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I455_Y_0 (.A(
        \sumreg[37]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I455_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I255_Y (.A(N740), .B(N732), .Y(
        N814));
    AO1 next_ireg_3_0_ADD_22x22_fast_I82_Y (.A(N355), .B(N352), .C(
        N351), .Y(N390));
    NOR2A inf_abs2_a_0_I_25 (.A(\DWACT_FINC_E_0[4] ), .B(integral[14]), 
        .Y(N_18));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I183_Y (.A(N659), .B(N655), .Y(
        N736));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I254_un1_Y (.A(N739), .B(N732), 
        .Y(I254_un1_Y));
    DFN1E1C0 \ireg[8]  (.D(\next_ireg_3[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[8]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I302_un1_Y (.A(N805), .B(N790), 
        .Y(I302_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I360_un1_Y (.A(N882), .B(N666), 
        .Y(I360_un1_Y));
    OA1 next_ireg_3_0_ADD_22x22_fast_I25_Y (.A(\i_adj[18]_net_1 ), .B(
        \i_adj[16]_net_1 ), .C(N312), .Y(N330));
    OA1 next_ireg_3_0_ADD_22x22_fast_I43_Y (.A(\i_adj[8]_net_1 ), .B(
        \i_adj[6]_net_1 ), .C(N288), .Y(N348));
    XNOR2 inf_abs1_a_2_I_35 (.A(sr_new[12]), .B(N_2), .Y(
        \inf_abs1_a_2[12] ));
    DFN1E1C0 \preg[8]  (.D(\p_adj[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[8]_net_1 ));
    XA1 \ireg_RNIURNG[23]  (.A(integral_1_0), .B(\ireg[23]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[23] ));
    XNOR2 inf_abs2_a_0_I_53 (.A(integral[24]), .B(N_9_0), .Y(
        \inf_abs2_a_0[18] ));
    DFN1E1C0 \i_adj[14]  (.D(\inf_abs2_5[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[14]_net_1 ));
    DFN1E1C0 \sumreg[32]  (.D(\next_sum[32] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[32]_net_1 ));
    XA1 \ireg_RNIE6AJ[5]  (.A(integral_1_0), .B(\ireg[5]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[5] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I346_Y (.A(
        ADD_40x40_fast_I346_un1_Y_0), .B(N1085), .C(
        ADD_40x40_fast_I346_Y_0), .Y(N1037));
    AO1 next_ireg_3_0_ADD_22x22_fast_I28_Y (.A(N305), .B(N309), .C(
        N308), .Y(N333));
    NOR3A un1_sumreg_0_0_ADD_40x40_fast_I25_G0N (.A(\sumreg[25]_net_1 )
        , .B(\ireg_m[25] ), .C(\un1_next_sum_0_iv_1[25] ), .Y(N546));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I249_Y (.A(N734), .B(N726), .Y(
        N808));
    NOR3B \ireg_RNIQMMG[10]  (.A(integral_1_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[10]_net_1 ), .Y(\un3_next_sum_m[10] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I351_Y (.A(
        ADD_40x40_fast_I351_un1_Y_0), .B(N1100), .C(
        ADD_40x40_fast_I351_Y_0), .Y(N1052));
    MX2 \i_adj_RNO[6]  (.A(integral[12]), .B(\inf_abs2_a_0[6] ), .S(
        integral_0_0), .Y(\inf_abs2_5[6] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I188_Y (.A(N664), .B(N661), .C(
        N660), .Y(N741));
    AND3 inf_abs1_a_2_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(N_6_0));
    OR2 \ireg_RNIDJQ41[20]  (.A(\un1_next_sum_iv_0[20] ), .B(
        \un1_next_sum_2[4] ), .Y(\un1_next_sum[20] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I17_P0N (.A(
        \un1_next_sum_iv_1[17] ), .B(\un1_next_sum_iv_2[17] ), .C(
        sum_17), .Y(N523));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I16_P0N (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(N520));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I49_Y (.A(\sumreg[33]_net_1 ), 
        .B(\sumreg[34]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N599)
        );
    XNOR2 inf_abs2_a_0_I_26 (.A(integral[15]), .B(N_18), .Y(
        \inf_abs2_a_0[9] ));
    NOR2A \sumreg_RNO[12]  (.A(\un1_sumreg[12] ), .B(\state[2]_net_1 ), 
        .Y(\next_sum[12] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I54_Y (.A(\sumreg[30]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N604)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I315_Y (.A(N804), .B(N819), .C(
        N803), .Y(N1088));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I112_Y (.A(sum_1_d0), .B(
        sum_2_d0), .C(\un1_next_sum[0] ), .Y(N662));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I177_Y_0 (.A(\i_adj[19]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(ADD_22x22_fast_I177_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I106_Y (.A(N483), .B(N487), .C(
        N486), .Y(N656));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I7_G0N (.A(\un1_next_sum[7] ), 
        .B(sum_7), .Y(N492_0));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I164_Y (.A(\i_adj[4]_net_1 ), .B(
        \i_adj[6]_net_1 ), .C(N394), .Y(\next_ireg_3[10] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_1 (.A(
        ADD_22x22_fast_I142_Y_0_a3_0), .B(N329), .C(
        ADD_22x22_fast_I142_Y_0_0), .Y(ADD_22x22_fast_I142_Y_0_1));
    XNOR2 inf_abs2_a_0_I_62 (.A(integral[25]), .B(N_6), .Y(
        \inf_abs2_a_0[21] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I419_Y_0 (.A(sum_1_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I419_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I68_Y (.A(N540), .B(N544), .C(
        N543), .Y(N618));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I22_G0N (.A(\un1_next_sum_2[4] ), 
        .B(\un1_next_sum_iv_0[22] ), .C(sum_22), .Y(N537));
    NOR2 inf_abs2_a_0_I_38 (.A(integral[18]), .B(integral[19]), .Y(
        \DWACT_FINC_E[8] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I380_Y_2 (.A(N758), .B(N773), .C(
        ADD_40x40_fast_I380_Y_1), .Y(ADD_40x40_fast_I380_Y_2));
    NOR3 inf_abs2_a_0_I_41 (.A(integral[19]), .B(integral[18]), .C(
        integral[20]), .Y(\DWACT_FINC_E[9] ));
    MX2 \p_adj_RNO[9]  (.A(sr_new[9]), .B(\inf_abs1_a_2[9] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[9] ));
    DFN1E1C0 \sumreg[33]  (.D(\next_sum[33] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[33]_net_1 ));
    XA1B \sumreg_RNO[2]  (.A(N745), .B(ADD_40x40_fast_I420_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[2] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I156_Y (.A(N632), .B(N629), .C(
        N628), .Y(N709));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I352_un1_Y_0 (.A(N798), .B(
        N782), .Y(ADD_40x40_fast_I352_un1_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I100_Y (.A(N492_0), .B(N496), .C(
        N495), .Y(N650));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I165_Y_0 (.A(\i_adj[7]_net_1 ), 
        .B(\i_adj[5]_net_1 ), .Y(ADD_22x22_fast_I165_Y_0));
    DFN1E1C0 \i_adj[12]  (.D(\inf_abs2_5[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[12]_net_1 ));
    AO1 \ireg_RNIJPU91[15]  (.A(\ireg[15]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[15] ), .Y(
        \un1_next_sum_iv_1[15] ));
    NOR2B \i_adj_RNO[19]  (.A(\inf_abs2_a_0[19] ), .B(integral[25]), 
        .Y(\inf_abs2_5[19] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I359_un1_Y (.A(N796), .B(N812), 
        .C(N745), .Y(I359_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I39_Y (.A(N291), .B(N294), .Y(
        N344));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I143_un1_Y_0 (.A(N375), .B(N367)
        , .C(N359), .Y(ADD_22x22_fast_I143_un1_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y_0 (.A(N335), .B(N332), .C(
        N331), .Y(ADD_22x22_fast_I126_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I14_G0N (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .Y(N308));
    DFN1E1C0 \sumreg[30]  (.D(\next_sum[30] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[30]_net_1 ));
    AND3 inf_abs2_a_0_I_39 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E_0[7] ), .C(\DWACT_FINC_E[8] ), .Y(N_13));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I24_Y (.A(N311), .B(
        \i_adj[18]_net_1 ), .C(\i_adj[16]_net_1 ), .Y(N329));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I37_Y (.A(N294), .B(N297), .Y(
        N342));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I302_Y (.A(I302_un1_Y), .B(N789), 
        .Y(N873));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I130_Y (.A(N606), .B(N602), .Y(
        N683));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I80_Y (.A(N522_0), .B(N526), .C(
        N525_0), .Y(N630));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I346_un1_Y_0 (.A(N786), .B(
        N770), .Y(ADD_40x40_fast_I346_un1_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I288_un1_Y (.A(N791), .B(N776), 
        .Y(I288_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I0_G0N (.A(N_228), .B(sum_0_d0)
        , .Y(N471));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I150_Y (.A(N626), .B(N623), .C(
        N622), .Y(N703));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I161_Y (.A(N637), .B(N633), .Y(
        N714));
    AO1 next_ireg_3_0_ADD_22x22_fast_I40_Y (.A(N287), .B(N291), .C(
        N290), .Y(N345));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I172_Y_0 (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[12]_net_1 ), .Y(ADD_22x22_fast_I172_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I346_Y_0 (.A(N785), .B(N770), .C(
        N769), .Y(ADD_40x40_fast_I346_Y_0));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I63_Y (.A(\sumreg[26]_net_1 ), 
        .B(\sumreg[27]_net_1 ), .C(\un1_next_sum_1_iv[26] ), .Y(N613));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I187_Y (.A(
        ADD_40x40_fast_I187_Y_0), .B(N659), .Y(N740));
    XA1B \sumreg_RNO[4]  (.A(N823), .B(ADD_40x40_fast_I422_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I352_Y (.A(
        ADD_40x40_fast_I352_un1_Y_0), .B(N1103), .C(
        ADD_40x40_fast_I352_Y_0), .Y(N1055));
    XA1B \sumreg_RNO[5]  (.A(N821), .B(ADD_40x40_fast_I423_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[5] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I378_Y (.A(N869), .B(N838), .C(
        ADD_40x40_fast_I378_Y_4), .Y(N1021));
    OR3 \ireg_RNICQ2H1[14]  (.A(\un24_next_sum_m[14] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[14] ), .Y(
        \un1_next_sum_iv_2[14] ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I45_Y (.A(\i_adj[8]_net_1 ), .B(
        \i_adj[6]_net_1 ), .C(N282), .Y(N350));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I171_Y (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .C(N513), .Y(\next_ireg_3[17] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_0_o3_0_0 (.A(N337), .B(
        N334), .C(N333), .Y(ADD_22x22_fast_I142_Y_0_o3_0_0));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I432_Y_0 (.A(
        \un1_next_sum_iv_1[14] ), .B(\un1_next_sum_iv_2[14] ), .C(
        sum_14), .Y(ADD_40x40_fast_I432_Y_0));
    DFN1E1C0 \sumreg[37]  (.D(\next_sum[37] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[37]_net_1 ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I51_Y (.A(\sumreg[32]_net_1 ), 
        .B(\sumreg[33]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N601)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I383_Y_1 (.A(N764), .B(N779), .C(
        ADD_40x40_fast_I383_Y_0), .Y(ADD_40x40_fast_I383_Y_1));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I23_P0N (.A(\un1_next_sum[23] ), 
        .B(sum_23), .Y(N541));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_2 (.A(N367), .B(N374), .C(
        ADD_22x22_fast_I143_Y_1), .Y(ADD_22x22_fast_I143_Y_2));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I66_Y (.A(N543), .B(N547), .C(
        N546), .Y(N616));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I445_Y_0 (.A(
        \sumreg[27]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I445_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I298_un1_Y (.A(N801), .B(N786), 
        .Y(I298_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I109_Y (.A(N481), .B(N484), .Y(
        N659));
    XNOR2 inf_abs2_a_0_I_28 (.A(integral[16]), .B(N_17), .Y(
        \inf_abs2_a_0[10] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I19_P0N (.A(\un1_next_sum[19] ), 
        .B(sum_19), .Y(N529));
    NOR3 inf_abs2_a_0_I_33 (.A(integral[17]), .B(integral[16]), .C(
        integral[15]), .Y(\DWACT_FINC_E_0[7] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I55_Y (.A(\sumreg[30]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N605)
        );
    DFN1C0 \state_1[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_1[2]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I48_Y (.A(N275), .B(N279), .C(
        N278), .Y(N353));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I3_G0N (.A(sum_3), .B(
        \un1_next_sum[0] ), .Y(N480));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I344_un1_Y (.A(N852), .B(N883), 
        .Y(I344_un1_Y));
    MX2 \i_adj_RNO[4]  (.A(integral[10]), .B(\inf_abs2_a_0[4] ), .S(
        integral_0_0), .Y(\inf_abs2_5[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I210_Y (.A(N695), .B(N688), .C(
        N687), .Y(N769));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I15_G0N (.A(
        \un1_next_sum_iv_1[15] ), .B(\un1_next_sum_iv_2[15] ), .C(
        sum_15), .Y(N516));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I425_Y_0 (.A(sum_7), .B(
        \un1_next_sum[7] ), .Y(ADD_40x40_fast_I425_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I139_Y (.A(N611), .B(N615), .Y(
        N692));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I384_un1_Y (.A(N882), .B(N666), 
        .C(N850), .Y(I384_un1_Y));
    NOR3B \preg_RNI3JN01[15]  (.A(sr_new_1_0), .B(\state[5]_net_1 ), 
        .C(\preg[15]_net_1 ), .Y(\un24_next_sum_m[15] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I277_Y (.A(N764), .B(N780), .Y(
        N848));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I159_Y (.A(N635), .B(N631), .Y(
        N712));
    DFN1E1C0 \i_adj[13]  (.D(\inf_abs2_5[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[13]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I104_Y (.A(N486), .B(N490), .C(
        N489), .Y(N654));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I115_un1_Y (.A(N393), .B(N266), 
        .Y(I115_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I54_un1_Y (.A(N270), .B(N266), 
        .Y(I54_un1_Y));
    NOR3 inf_abs2_a_0_I_29 (.A(integral[13]), .B(integral[12]), .C(
        integral[14]), .Y(\DWACT_FINC_E[5] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I130_Y_0 (.A(N386), .B(N379), .C(
        N378), .Y(ADD_22x22_fast_I130_Y_0));
    DFN1E1C0 \preg[12]  (.D(\p_adj[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[12]_net_1 ));
    MX2 \i_adj_RNO[2]  (.A(integral[8]), .B(\inf_abs2_a_0[2] ), .S(
        integral_0_0), .Y(\inf_abs2_5[2] ));
    DFN1E1C0 \i_adj[5]  (.D(\inf_abs2_5[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[5]_net_1 ));
    DFN1E1C0 \ireg[20]  (.D(\next_ireg_3[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[20]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I379_Y_0 (.A(\sumreg[37]_net_1 )
        , .B(\sumreg[36]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(
        ADD_40x40_fast_I379_Y_0));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I321_un1_Y (.A(N734), .B(
        ADD_40x40_fast_I257_Y_1), .C(\un1_next_sum[0] ), .Y(I321_un1_Y)
        );
    OR3 un1_sumreg_0_0_ADD_m8_i_o4_1 (.A(sum_2_d0), .B(sum_1_d0), .C(
        sum_0_d0), .Y(ADD_m8_i_o4_1));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I378_Y_0 (.A(\sumreg[38]_net_1 )
        , .B(\sumreg[37]_net_1 ), .C(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I378_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I134_Y (.A(N610), .B(N606), .Y(
        N687));
    DFN1E1C0 \i_adj[0]  (.D(\inf_abs2_5[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[0]_net_1 ));
    DFN1E1C0 \p_adj[6]  (.D(\inf_abs1_5[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[6]_net_1 ));
    MX2 \p_adj_RNO[4]  (.A(sr_new[4]), .B(\inf_abs1_a_2[4] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I154_Y (.A(N630), .B(N627), .C(
        N626), .Y(N707));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I211_Y (.A(N688), .B(N696), .Y(
        N770));
    OR3 \ireg_RNIGU2H1[16]  (.A(\un24_next_sum_m[16] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[16] ), .Y(
        \un1_next_sum_iv_2[16] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I12_G0N (.A(
        \un1_next_sum_iv_1[12] ), .B(\un1_next_sum_iv_2[12] ), .C(
        sum_12), .Y(N507_0));
    XA1B \sumreg_RNO[24]  (.A(N1058), .B(ADD_40x40_fast_I442_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[24] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I59_Y (.A(N328), .B(N332), .Y(
        N367));
    MX2 \i_adj_RNO[0]  (.A(integral[6]), .B(integral[6]), .S(
        integral_0_0), .Y(\inf_abs2_5[0] ));
    AND3 inf_abs2_a_0_I_42 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E_0[7] ), .C(\DWACT_FINC_E[9] ), .Y(N_12_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I17_P0N_i_o3 (.A(
        \i_adj[19]_net_1 ), .B(\i_adj[17]_net_1 ), .Y(N_9));
    OR2 \ireg_RNI0O333[11]  (.A(\un1_next_sum_iv_2[11] ), .B(
        \un1_next_sum_iv_1[11] ), .Y(\un1_next_sum[11] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I218_Y (.A(N703), .B(N696), .C(
        N695), .Y(N777));
    XNOR2 inf_abs2_a_0_I_23 (.A(integral[14]), .B(N_19), .Y(
        \inf_abs2_a_0[8] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I66_Y (.A(N339), .B(N336), .C(
        N335), .Y(N374));
    XA1 \ireg_RNID5AJ[4]  (.A(integral_1_0), .B(\ireg[4]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[4] ));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I44_Y (.A(N281), .B(
        \i_adj[8]_net_1 ), .C(\i_adj[6]_net_1 ), .Y(N349));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I439_Y_0 (.A(sum_21), .B(
        \un1_next_sum[21] ), .Y(ADD_40x40_fast_I439_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I450_Y_0 (.A(
        \sumreg[32]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I450_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I234_Y (.A(N719), .B(N712), .C(
        N711), .Y(N793));
    NOR3 inf_abs1_a_2_I_33 (.A(sr_new[10]), .B(sr_new[9]), .C(
        sr_new[11]), .Y(\DWACT_FINC_E[7] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I384_Y (.A(I384_un1_Y), .B(
        ADD_40x40_fast_I384_Y_1), .C(I342_un1_Y), .Y(N1033));
    MX2 \i_adj_RNO[7]  (.A(integral[13]), .B(\inf_abs2_a_0[7] ), .S(
        integral_0_0), .Y(\inf_abs2_5[7] ));
    DFN1E1C0 \i_adj[21]  (.D(\inf_abs2_5[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[21]_net_1 ));
    XA1B \sumreg_RNO[9]  (.A(N1103), .B(ADD_40x40_fast_I427_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[9] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I59_Y (.A(\sumreg[29]_net_1 ), 
        .B(\sumreg[28]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N609)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I162_Y (.A(N638), .B(N635), .C(
        N634), .Y(N715));
    NOR3B \ireg_RNIJK7M_0[9]  (.A(\state[3]_net_1 ), .B(
        \ireg[9]_net_1 ), .C(integral[25]), .Y(\ireg_m[9] ));
    DFN1E1C0 \ireg[14]  (.D(\next_ireg_3[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[14]_net_1 ));
    DFN1E1C0 \p_adj[11]  (.D(\inf_abs1_5[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[11]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I82_Y (.A(N519), .B(N523), .C(
        N522_0), .Y(N632));
    DFN1E1C0 \i_adj[16]  (.D(\inf_abs2_5[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[16]_net_1 ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I4_P0N (.A(\i_adj[4]_net_1 ), .B(
        \i_adj[6]_net_1 ), .Y(N279));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I178_Y_0 (.A(\i_adj[20]_net_1 ), 
        .B(\i_adj[18]_net_1 ), .Y(ADD_22x22_fast_I178_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I131_Y_0 (.A(N345), .B(N342), .C(
        N341), .Y(ADD_22x22_fast_I131_Y_0));
    NOR3B \ireg_RNIJK7M[9]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[9]_net_1 ), .Y(\un3_next_sum_m[9] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I437_Y_0 (.A(sum_19), .B(
        \un1_next_sum[19] ), .Y(ADD_40x40_fast_I437_Y_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I13_P0N (.A(
        \un1_next_sum_iv_1[13] ), .B(\un1_next_sum_iv_2[13] ), .C(
        sum_13), .Y(N511));
    AO1 next_ireg_3_0_ADD_22x22_fast_I32_Y (.A(N299), .B(N303), .C(
        N302), .Y(N337));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I352_Y_0 (.A(N797), .B(N782), .C(
        N781), .Y(ADD_40x40_fast_I352_Y_0));
    MX2 \i_adj_RNO[11]  (.A(integral[17]), .B(\inf_abs2_a_0[11] ), .S(
        integral_0_0), .Y(\inf_abs2_5[11] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I15_G0N (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(N311));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I298_Y (.A(I298_un1_Y), .B(N785), 
        .Y(N869));
    DFN1E1C0 \ireg[4]  (.D(\i_adj[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[4]_net_1 ));
    OR2 \preg_RNIGMHS[9]  (.A(next_sum_0_sqmuxa_1), .B(
        \un24_next_sum_m[9] ), .Y(\un1_next_sum_iv_0[9] ));
    MX2 \p_adj_RNO[11]  (.A(sr_new[11]), .B(\inf_abs1_a_2[11] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[11] ));
    AX1D next_ireg_3_0_ADD_22x22_fast_I172_Y (.A(I130_un1_Y), .B(
        ADD_22x22_fast_I130_Y_0), .C(ADD_22x22_fast_I172_Y_0), .Y(
        \next_ireg_3[18] ));
    XA1B \sumreg_RNO[37]  (.A(N1025), .B(ADD_40x40_fast_I455_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[37] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I381_un1_Y (.A(N876), .B(N823), 
        .C(N844), .Y(I381_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I141_Y (.A(N613), .B(N617), .Y(
        N694));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I83_Y (.A(N356), .B(N352), .Y(
        N391));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I111_Y (.A(N393), .B(N385), .Y(
        N425));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I175_Y (.A(N647), .B(N651), .Y(
        N728));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I378_un1_Y_0 (.A(N786), .B(
        N802), .C(N817), .Y(ADD_40x40_fast_I378_un1_Y_0));
    DFN1E1C0 \sumreg[24]  (.D(\next_sum[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(\sumreg[24]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I26_Y (.A(N308), .B(N312), .C(
        N311), .Y(N331));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I24_G0N (.A(\un1_next_sum[24] )
        , .B(\sumreg[24]_net_1 ), .Y(N543));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I175_Y (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .C(N_11), .Y(\next_ireg_3[21] ));
    NOR3B \ireg_RNIJCK8[18]  (.A(integral_1_0), .B(\state[3]_net_1 ), 
        .C(\ireg[18]_net_1 ), .Y(\un3_next_sum_m[18] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I431_Y_0 (.A(
        \un1_next_sum_iv_1[13] ), .B(\un1_next_sum_iv_2[13] ), .C(
        sum_13), .Y(ADD_40x40_fast_I431_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I300_Y (.A(I300_un1_Y), .B(N787), 
        .Y(N871));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I382_un1_Y_0 (.A(N743), .B(
        N878), .Y(ADD_40x40_fast_I382_un1_Y_0));
    NOR2B \state_RNIBU9J[3]  (.A(\state[3]_net_1 ), .B(integral[25]), 
        .Y(next_sum_0_sqmuxa));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I103_Y (.A(N490), .B(N493), .Y(
        N653));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I88_Y (.A(N510), .B(N514), .C(
        N513_0), .Y(N638));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I0_P0N (.A(N_228), .B(sum_0_d0), 
        .Y(N472));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I260_Y (.A(N740), .B(N666), .C(
        N739), .Y(N821));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I8_P0N (.A(
        \un1_next_sum_iv_1[8] ), .B(\un1_next_sum_iv_2[8] ), .C(sum_8), 
        .Y(N496));
    OR3 \state_RNITOC71[4]  (.A(next_sum_1_sqmuxa_2), .B(
        next_sum_1_sqmuxa_1), .C(next_sum_1_sqmuxa), .Y(
        \un1_next_sum_1_iv_0[26] ));
    OR2 \ireg_RNIGMQ41[23]  (.A(\un1_next_sum_iv_0[23] ), .B(
        \un1_next_sum_2[4] ), .Y(\un1_next_sum[23] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I216_un1_Y (.A(N701), .B(N694), 
        .Y(I216_un1_Y));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I379_un1_Y_0 (.A(N788), .B(
        N804), .C(N840), .Y(ADD_40x40_fast_I379_un1_Y_0));
    NOR2B \state_RNIAMDD[0]  (.A(sum_enable), .B(sum_rdy), .Y(
        \state_RNIAMDD[0]_net_1 ));
    MX2 \i_adj_RNO[15]  (.A(integral[21]), .B(\inf_abs2_a_0[15] ), .S(
        integral_0_0), .Y(\inf_abs2_5[15] ));
    DFN1E1C0 \sumreg[14]  (.D(\next_sum[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_14));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I350_Y (.A(I290_un1_Y), .B(N777), 
        .C(I350_un1_Y), .Y(N1049));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I203_Y (.A(N680), .B(N688), .Y(
        N762));
    NOR2B \i_adj_RNO[20]  (.A(\inf_abs2_a_0[20] ), .B(integral[25]), 
        .Y(\inf_abs2_5[20] ));
    XNOR2 inf_abs1_a_2_I_14 (.A(sr_new[5]), .B(N_9_1), .Y(
        \inf_abs1_a_2[5] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I170_Y_0 (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[12]_net_1 ), .Y(ADD_22x22_fast_I170_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I133_Y (.A(N605), .B(N609), .Y(
        N686));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I215_Y (.A(N700), .B(N692), .Y(
        N774));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I279_Y (.A(N766), .B(N782), .Y(
        N850));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I153_Y (.A(N625), .B(N629), .Y(
        N706));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I79_Y (.A(N348), .B(N352), .Y(
        N387));
    XA1B \sumreg_RNO[30]  (.A(N1040), .B(ADD_40x40_fast_I448_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[30] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I77_Y (.A(N350), .B(N346), .Y(
        N385));
    OR3 \ireg_RNIK23H1[18]  (.A(\un24_next_sum_m[18] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[18] ), .Y(
        \un1_next_sum_iv_2[18] ));
    XNOR2 inf_abs2_a_0_I_9 (.A(integral[9]), .B(N_24), .Y(
        \inf_abs2_a_0[3] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I233_Y (.A(N641), .B(N637), .C(
        N710), .Y(N792));
    XA1B \sumreg_RNO[31]  (.A(N1037), .B(ADD_40x40_fast_I449_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[31] ));
    NOR3 inf_abs2_a_0_I_10 (.A(integral[7]), .B(integral[6]), .C(
        integral[8]), .Y(\DWACT_FINC_E_0[0] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I440_Y_0 (.A(
        \un1_next_sum_2[4] ), .B(\un1_next_sum_iv_0[22] ), .C(sum_22), 
        .Y(ADD_40x40_fast_I440_Y_0));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I253_Y (.A(N653), .B(N649), .C(
        N738), .Y(N812));
    OR3 \preg_RNI19PI1[8]  (.A(\un24_next_sum_m[8] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[8] ), .Y(
        \un1_next_sum_iv_2[8] ));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I52_Y (.A(N269), .B(
        \i_adj[4]_net_1 ), .C(\i_adj[2]_net_1 ), .Y(N357));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I108_Y (.A(N480), .B(N484), .C(
        N483), .Y(N658));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I261_Y (.A(I116_un1_Y), .B(N741), 
        .Y(N823));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I173_Y (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[15]_net_1 ), .C(N507), .Y(\next_ireg_3[19] ));
    NOR2 inf_abs1_a_2_I_15 (.A(sr_new[3]), .B(sr_new[4]), .Y(
        \DWACT_FINC_E_0[1] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I83_Y (.A(N520), .B(N523), .Y(
        N633));
    XA1B \sumreg_RNO[25]  (.A(N1055), .B(ADD_40x40_fast_I443_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[25] ));
    DFN1E1C0 \i_adj[11]  (.D(\inf_abs2_5[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[11]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I307_Y (.A(N810), .B(N794), .Y(
        N878));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I138_Y (.A(N614), .B(N611), .C(
        N610), .Y(N691));
    DFN1E1C0 \ireg[11]  (.D(\next_ireg_3[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[11]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I311_Y (.A(N814), .B(N798), .Y(
        N882));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I420_Y_0 (.A(sum_2_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I420_Y_0));
    DFN1C0 \state[3]  (.D(\state[6]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[3]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I158_Y (.A(N634), .B(N631), .C(
        N630), .Y(N711));
    MX2 \i_adj_RNO[17]  (.A(integral[23]), .B(\inf_abs2_a_0[17] ), .S(
        integral_0_0), .Y(\inf_abs2_5[17] ));
    DFN1E1C0 \i_adj[1]  (.D(\inf_abs2_5[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[1]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I80_Y (.A(N353), .B(N350), .C(
        N349), .Y(N388));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I86_Y (.A(N513_0), .B(N517), .C(
        N516), .Y(N636));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I236_Y (.A(N721), .B(N714), .C(
        N713), .Y(N795));
    DFN1E1C0 \sumreg[3]  (.D(\next_sum[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_3));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I358_un1_Y (.A(N878), .B(N743), 
        .Y(I358_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I220_Y (.A(N705), .B(N698), .C(
        N697), .Y(N779));
    DFN1E1C0 \sumreg_1[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(sum_1_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I382_Y_1 (.A(N762), .B(N777), .C(
        ADD_40x40_fast_I382_Y_0), .Y(ADD_40x40_fast_I382_Y_1));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I4_G0N (.A(\i_adj[4]_net_1 ), 
        .B(\i_adj[6]_net_1 ), .Y(N278));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I357_Y (.A(N876), .B(N823), .C(
        N875), .Y(N1070));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I85_Y (.A(
        ADD_22x22_fast_I85_Y_0), .B(N354), .Y(N393));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I24_P0N (.A(\un1_next_sum[24] ), 
        .B(\sumreg[24]_net_1 ), .Y(N544));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I142_Y (.A(N618), .B(N615), .C(
        N614), .Y(N695));
    OR3 \ireg_RNIES2H1[15]  (.A(\un24_next_sum_m[15] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[15] ), .Y(
        \un1_next_sum_iv_2[15] ));
    DFN1C0 \state_0[1]  (.D(\state_RNIAMDD[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_0[1]_net_1 ));
    NOR3 inf_abs2_a_0_I_50 (.A(integral[22]), .B(integral[21]), .C(
        integral[23]), .Y(\DWACT_FINC_E[12] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I347_un1_Y_0 (.A(N788), .B(
        N772), .Y(ADD_40x40_fast_I347_un1_Y_0));
    NOR3B \ireg_RNIIBK8[17]  (.A(integral_1_0), .B(\state[3]_net_1 ), 
        .C(\ireg[17]_net_1 ), .Y(\un3_next_sum_m[17] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I3_G0N (.A(\i_adj[3]_net_1 ), 
        .B(\i_adj[5]_net_1 ), .Y(N275));
    XNOR2 inf_abs1_a_2_I_9 (.A(sr_new[3]), .B(N_11_1), .Y(
        \inf_abs1_a_2[3] ));
    NOR3B inf_abs1_a_2_I_16 (.A(\DWACT_FINC_E_0[1] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[5]), .Y(N_8_0));
    NOR2B \preg_RNIIIAM[14]  (.A(\preg[14]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[14] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I355_un1_Y (.A(N788), .B(N804), 
        .C(N819), .Y(I355_un1_Y));
    AO1 next_ireg_3_0_ADD_22x22_fast_I46_Y (.A(N278), .B(N282), .C(
        N281), .Y(N351));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I13_G0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[15]_net_1 ), .Y(N305));
    AO1 \ireg_RNINTU91[17]  (.A(\ireg[17]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[17] ), .Y(
        \un1_next_sum_iv_1[17] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I361_un1_Y (.A(N884), .B(
        \un1_next_sum[0] ), .Y(I361_un1_Y));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I350_un1_Y (.A(N778), .B(N794), 
        .C(N1097), .Y(I350_un1_Y));
    VCC VCC_i (.Y(VCC));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I221_Y (.A(N698), .B(N706), .Y(
        N780));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I14_G0N (.A(
        \un1_next_sum_iv_1[14] ), .B(\un1_next_sum_iv_2[14] ), .C(
        sum_14), .Y(N513_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I116_Y (.A(I116_un1_Y), .B(N471), 
        .Y(N666));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I50_Y (.A(\sumreg[33]_net_1 ), 
        .B(\sumreg[32]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N600)
        );
    AND3 inf_abs1_a_2_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(
        \DWACT_FINC_E[4] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I6_G0N (.A(\un1_next_sum[6] ), 
        .B(sum_6), .Y(N489));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I385_Y_1 (.A(I208_un1_Y), .B(
        N685), .C(I280_un1_Y), .Y(ADD_40x40_fast_I385_Y_1));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I383_un1_Y (.A(
        ADD_40x40_fast_I383_un1_Y_0), .B(N848), .Y(I383_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I185_Y (.A(N661), .B(N657), .Y(
        N738));
    OA1 next_ireg_3_0_ADD_22x22_fast_I85_Y_0 (.A(\i_adj[4]_net_1 ), .B(
        \i_adj[2]_net_1 ), .C(N270), .Y(ADD_22x22_fast_I85_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I448_Y_0 (.A(
        \sumreg[30]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I448_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I107_Y (.A(N484), .B(N487), .Y(
        N657));
    AO1 next_ireg_3_0_ADD_22x22_fast_I129_Y_0 (.A(N384), .B(N377), .C(
        N376), .Y(ADD_22x22_fast_I129_Y_0));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I130_un1_Y (.A(N379), .B(N387), 
        .C(N394), .Y(I130_un1_Y));
    AO1 next_ireg_3_0_ADD_22x22_fast_I112_Y (.A(N387), .B(N394), .C(
        N386), .Y(N522));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I228_Y (.A(N713), .B(N706), .C(
        N705), .Y(N787));
    NOR3 inf_abs1_a_2_I_8 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2]), 
        .Y(N_11_1));
    XA1B \sumreg_RNO[26]  (.A(N1052), .B(ADD_40x40_fast_I444_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[26] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I378_Y_4 (.A(
        ADD_40x40_fast_I378_un1_Y_0), .B(N838), .C(
        ADD_40x40_fast_I378_Y_3), .Y(ADD_40x40_fast_I378_Y_4));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I454_Y_0 (.A(
        \sumreg[36]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I454_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I110_Y (.A(sum_2_d0), .B(
        \un1_next_sum[0] ), .C(N480), .Y(N660));
    XA1B \sumreg_RNO[17]  (.A(N1079), .B(ADD_40x40_fast_I435_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[17] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I359_Y (.A(N795), .B(I308_un1_Y), 
        .C(I359_un1_Y), .Y(N1076));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I137_Y (.A(N613), .B(N609), .Y(
        N690));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I129_un1_Y_0 (.A(N385), .B(N377)
        , .Y(ADD_22x22_fast_I129_un1_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I453_Y_0 (.A(
        \sumreg[35]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I453_Y_0));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I48_Y (.A(\sumreg[33]_net_1 ), 
        .B(\sumreg[34]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(
        I122_un1_Y));
    NOR2A inf_abs1_a_2_I_25 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .Y(
        N_5));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I157_Y (.A(N633), .B(N629), .Y(
        N710));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I428_Y_0 (.A(
        \un1_next_sum_iv_1[10] ), .B(\un1_next_sum_iv_2[10] ), .C(
        sum_10), .Y(ADD_40x40_fast_I428_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I312_Y (.A(I312_un1_Y), .B(N799), 
        .Y(N883));
    DFN1E1C0 \preg[11]  (.D(\p_adj[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[11]_net_1 ));
    XA1B \sumreg_RNO[23]  (.A(N1061), .B(ADD_40x40_fast_I441_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[23] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I131_un1_Y (.A(
        ADD_22x22_fast_I131_un1_Y_0), .B(N396), .Y(I131_un1_Y));
    DFN1E1C0 \sumreg[22]  (.D(\next_sum[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(sum_22));
    NOR2B \preg_RNIMMAM[18]  (.A(\preg[18]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[18] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I115_Y (.A(I115_un1_Y), .B(N392), 
        .Y(N531));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I5_P0N (.A(\un1_next_sum[5] ), 
        .B(sum_5), .Y(N487));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I20_G0N (.A(\un1_next_sum[20] )
        , .B(sum_20), .Y(N531_0));
    DFN1E1C0 \ireg[13]  (.D(\next_ireg_3[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[13]_net_1 ));
    XA1B \sumreg_RNO[29]  (.A(N1043), .B(ADD_40x40_fast_I447_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[29] ));
    DFN1E1C0 \p_adj[8]  (.D(\inf_abs1_5[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[8]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I61_Y (.A(N334), .B(N330), .Y(
        N369));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I351_Y_0 (.A(N795), .B(N780), .C(
        N779), .Y(ADD_40x40_fast_I351_Y_0));
    AX1D next_ireg_3_0_ADD_22x22_fast_I177_Y (.A(I124_un1_Y), .B(
        ADD_22x22_fast_I144_Y_2), .C(ADD_22x22_fast_I177_Y_0), .Y(
        \next_ireg_3[23] ));
    OR2 \ireg_RNID8P71[6]  (.A(\un3_next_sum_m[6] ), .B(
        \un1_next_sum_iv_0[6] ), .Y(\un1_next_sum_iv_2[6] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I84_Y (.A(N357), .B(N354), .C(
        N353), .Y(N392));
    NOR3B \ireg_RNITPMG[13]  (.A(integral_1_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[13]_net_1 ), .Y(\un3_next_sum_m[13] ));
    NOR3B \ireg_RNIRNMG[11]  (.A(integral_1_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[11]_net_1 ), .Y(\un3_next_sum_m[11] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I240_Y (.A(I240_un1_Y), .B(N717), 
        .Y(N799));
    XNOR2 inf_abs1_a_2_I_7 (.A(sr_new[2]), .B(N_12), .Y(
        \inf_abs1_a_2[2] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I240_un1_Y (.A(N641), .B(N637), 
        .C(N725), .Y(I240_un1_Y));
    XNOR2 inf_abs2_a_0_I_17 (.A(integral[12]), .B(N_21), .Y(
        \inf_abs2_a_0[6] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I142_Y_0_a3_1_1 (.A(
        \i_adj[19]_net_1 ), .B(\i_adj[17]_net_1 ), .Y(N_14_1));
    DFN1E1C0 \sumreg[12]  (.D(\next_sum[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_12));
    DFN1E1C0 \ireg[15]  (.D(\next_ireg_3[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[15]_net_1 ));
    XA1B \sumreg_RNO[1]  (.A(N666), .B(ADD_40x40_fast_I419_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[1] ));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I179_Y (.A(\i_adj[19]_net_1 ), 
        .B(\i_adj[21]_net_1 ), .C(N492), .Y(\next_ireg_3[25] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I97_Y (.A(N499), .B(N502), .Y(
        N647));
    OR2 next_ireg_3_0_ADD_22x22_fast_I8_P0N (.A(\i_adj[10]_net_1 ), .B(
        \i_adj[8]_net_1 ), .Y(N291));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I280_un1_Y (.A(N694), .B(N686), 
        .C(N783), .Y(I280_un1_Y));
    DFN1E1C0 \sumreg_2[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNII1EM[6]_net_1 ), .Q(sum_2_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I7_P0N (.A(\i_adj[9]_net_1 ), .B(
        \i_adj[7]_net_1 ), .Y(N288));
    NOR3 inf_abs1_a_2_I_18 (.A(sr_new[4]), .B(sr_new[3]), .C(sr_new[5])
        , .Y(\DWACT_FINC_E_0[2] ));
    XNOR2 inf_abs1_a_2_I_26 (.A(sr_new[9]), .B(N_5), .Y(
        \inf_abs1_a_2[9] ));
    
endmodule


module sig_gen(
       vd_done,
       n_rst_c,
       clk_c,
       sig_old_i_0,
       sig_prev
    );
input  vd_done;
input  n_rst_c;
input  clk_c;
output sig_old_i_0;
output sig_prev;

    wire sig_prev_i, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(clk_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev_inst_1 (.D(vd_done), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(sig_prev));
    INV sig_old_RNO (.A(sig_prev), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module spi_stp_12s_1_1(
       cur_vd,
       N_29,
       din_12_c,
       n_rst_c,
       cur_clk
    );
output [11:0] cur_vd;
input  N_29;
input  din_12_c;
input  n_rst_c;
input  cur_clk;

    wire GND, VCC;
    
    DFN1E0C0 \sr[7]  (.D(cur_vd[6]), .CLK(cur_clk), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[7]));
    DFN1E0C0 \sr[5]  (.D(cur_vd[4]), .CLK(cur_clk), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[5]));
    DFN1E0C0 \sr[10]  (.D(cur_vd[9]), .CLK(cur_clk), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[10]));
    DFN1E0C0 \sr[8]  (.D(cur_vd[7]), .CLK(cur_clk), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[8]));
    DFN1E0C0 \sr[3]  (.D(cur_vd[2]), .CLK(cur_clk), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[3]));
    DFN1E0C0 \sr[1]  (.D(cur_vd[0]), .CLK(cur_clk), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[1]));
    DFN1E0C0 \sr[2]  (.D(cur_vd[1]), .CLK(cur_clk), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[2]));
    DFN1E0C0 \sr[9]  (.D(cur_vd[8]), .CLK(cur_clk), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[9]));
    VCC VCC_i (.Y(VCC));
    DFN1E0C0 \sr[11]  (.D(cur_vd[10]), .CLK(cur_clk), .CLR(n_rst_c), 
        .E(N_29), .Q(cur_vd[11]));
    DFN1E0C0 \sr[0]  (.D(din_12_c), .CLK(cur_clk), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[0]));
    GND GND_i (.Y(GND));
    DFN1E0C0 \sr[6]  (.D(cur_vd[5]), .CLK(cur_clk), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[6]));
    DFN1E0C0 \sr[4]  (.D(cur_vd[3]), .CLK(cur_clk), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[4]));
    
endmodule


module sig_gen_10_0(
       cs_i_1,
       n_rst_c,
       cur_clk,
       vd_done
    );
input  cs_i_1;
input  n_rst_c;
input  cur_clk;
output vd_done;

    wire sig_prev_i, sig_prev_net_1, sig_old_i_0, GND, VCC;
    
    NOR2B sig_old_RNI4485 (.A(sig_old_i_0), .B(sig_prev_net_1), .Y(
        vd_done));
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(cur_clk), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev (.D(cs_i_1), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        sig_prev_net_1));
    INV sig_old_RNO (.A(sig_prev_net_1), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module spi_ctl_12s_0(
       n_rst_c,
       cur_clk,
       N_29,
       cs_i_1,
       cs_i_1_i
    );
input  n_rst_c;
input  cur_clk;
output N_29;
output cs_i_1;
output cs_i_1_i;

    wire cnt_m1_0_a2_0, \cnt[14]_net_1 , \cnt[13]_net_1 , 
        cnt_m6_0_a2_6, cnt_m6_0_a2_0, \cnt[3]_net_1 , cnt_m5_0_a2_2, 
        cnt_m6_0_a2_2, \cnt[7]_net_1 , \cnt[8]_net_1 , \cnt[11]_net_1 , 
        \cnt[10]_net_1 , cnt_m7_0_a2_4, \cnt[5]_net_1 , cnt_m7_0_a2_3, 
        \cnt[6]_net_1 , cnt_m7_0_a2_1, \cnt[9]_net_1 , 
        state_tr0_0_a3_12, state_tr0_0_a3_6, state_tr0_0_a3_9, N_103, 
        \cnt[4]_net_1 , state_tr0_0_a3_8, state_tr0_0_a3_4, 
        state_tr0_0_a3_7, state_tr0_0_a3_2, \cnt[0]_net_1 , 
        \cnt[1]_net_1 , state_tr0_0_a3_1, \cnt[15]_net_1 , 
        \cnt[12]_net_1 , vd_stp_en_i_a3_9, vd_stp_en_i_a3_4, 
        vd_stp_en_i_a3_3, N_73, vd_stp_en_i_a3_8, vd_stp_en_i_a3_2, 
        vd_stp_en_i_a3_5, cnt_m6_0_a2_5_6, cnt_m6_0_a2_5_0, 
        cnt_m6_0_a2_5, \cnt[2]_net_1 , cnt_m5_0_a2_3, cnt_m2_0_a2_0, 
        cnt_m5_0_a2_1, cnt_m2_0_a2_2, cnt_m2_0_a2_1, N_74, 
        cnt_N_13_mux, N_33, N_31, cnt_N_7_mux_0_0, cnt_N_3_mux_0, 
        cnt_N_11_mux_2, cnt_N_15_mux, cnt_N_13_mux_0, N_30, 
        \state_RNO_0[0]_net_1 , N_26, N_24, N_22, N_20, N_97, N_18, 
        N_14, N_12, N_36, \cnt_RNO_2[6]_net_1 , cnt_n10, d_N_3_mux_3, 
        \cnt_RNO_1[10]_net_1 , cnt_n0, cnt_n15, cnt_n14, cnt_n13, N_72, 
        cnt_n12, cnt_n11, cnt_n9, N_38, GND, VCC;
    
    NOR2B \cnt_RNO_2[6]  (.A(\cnt[4]_net_1 ), .B(\cnt[3]_net_1 ), .Y(
        cnt_m2_0_a2_2));
    XA1A \cnt_RNO[8]  (.A(\cnt[8]_net_1 ), .B(N_36), .C(cs_i_1), .Y(
        N_12));
    NOR3C \cnt_RNO_3[10]  (.A(\cnt[3]_net_1 ), .B(\cnt[5]_net_1 ), .C(
        cs_i_1), .Y(cnt_m7_0_a2_4));
    NOR3A \state_RNO_0[0]  (.A(state_tr0_0_a3_4), .B(\cnt[6]_net_1 ), 
        .C(\cnt[7]_net_1 ), .Y(state_tr0_0_a3_8));
    NOR2 \cnt_RNI78RL[2]  (.A(\cnt[3]_net_1 ), .B(\cnt[2]_net_1 ), .Y(
        N_103));
    XA1A \cnt_RNO[2]  (.A(N_30), .B(\cnt[2]_net_1 ), .C(cs_i_1), .Y(
        N_24));
    NOR3C \cnt_RNI25NB1[9]  (.A(\cnt[9]_net_1 ), .B(\cnt[6]_net_1 ), 
        .C(cnt_m6_0_a2_2), .Y(cnt_m6_0_a2_5));
    DFN1C0 \cnt[2]  (.D(N_24), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[2]_net_1 ));
    NOR3B \cnt_RNISG6U3[3]  (.A(cnt_m6_0_a2_6), .B(cnt_m6_0_a2_5), .C(
        N_31), .Y(cnt_N_13_mux));
    NOR2 \cnt_RNIGHRL[6]  (.A(\cnt[8]_net_1 ), .B(\cnt[6]_net_1 ), .Y(
        vd_stp_en_i_a3_3));
    DFN1C0 \cnt[8]  (.D(N_12), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[8]_net_1 ));
    DFN1C0 \cnt[1]  (.D(N_26), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[1]_net_1 ));
    OA1C \cnt_RNO_0[4]  (.A(\cnt[3]_net_1 ), .B(N_31), .C(
        \cnt[4]_net_1 ), .Y(N_97));
    NOR3C \cnt_RNIHSMT1[10]  (.A(vd_stp_en_i_a3_2), .B(
        state_tr0_0_a3_1), .C(vd_stp_en_i_a3_5), .Y(vd_stp_en_i_a3_8));
    DFN1C0 \cnt[11]  (.D(cnt_n11), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[11]_net_1 ));
    NOR3C \cnt_RNO_0[6]  (.A(cnt_m2_0_a2_1), .B(cnt_m2_0_a2_0), .C(
        cnt_m2_0_a2_2), .Y(cnt_N_7_mux_0_0));
    NOR2B \cnt_RNO_1[15]  (.A(\cnt[14]_net_1 ), .B(\cnt[13]_net_1 ), 
        .Y(cnt_m1_0_a2_0));
    XA1A \cnt_RNO[3]  (.A(N_31), .B(\cnt[3]_net_1 ), .C(cs_i_1), .Y(
        N_22));
    OR2B \cnt_RNO_0[13]  (.A(cnt_N_13_mux), .B(\cnt[12]_net_1 ), .Y(
        N_72));
    NOR2B \cnt_RNIABRL[2]  (.A(\cnt[2]_net_1 ), .B(\cnt[6]_net_1 ), .Y(
        cnt_m5_0_a2_1));
    NOR3B \state_RNO_6[0]  (.A(\cnt[5]_net_1 ), .B(N_103), .C(
        \cnt[4]_net_1 ), .Y(state_tr0_0_a3_9));
    VCC VCC_i (.Y(VCC));
    XA1 \cnt_RNO[1]  (.A(\cnt[0]_net_1 ), .B(\cnt[1]_net_1 ), .C(
        cs_i_1), .Y(N_26));
    NOR2 \cnt_RNIIJRL[9]  (.A(\cnt[9]_net_1 ), .B(\cnt[7]_net_1 ), .Y(
        vd_stp_en_i_a3_4));
    NOR2B \cnt_RNIHIRL[7]  (.A(\cnt[7]_net_1 ), .B(\cnt[8]_net_1 ), .Y(
        cnt_m6_0_a2_2));
    OR2B \cnt_RNI49DN2[7]  (.A(cnt_N_11_mux_2), .B(\cnt[7]_net_1 ), .Y(
        N_36));
    DFN1C0 \cnt[6]  (.D(\cnt_RNO_2[6]_net_1 ), .CLK(cur_clk), .CLR(
        n_rst_c), .Q(\cnt[6]_net_1 ));
    NOR3C \cnt_RNO_0[15]  (.A(cnt_m1_0_a2_0), .B(\cnt[12]_net_1 ), .C(
        cnt_N_13_mux), .Y(cnt_N_3_mux_0));
    NOR2 \cnt_RNI8MTG[11]  (.A(\cnt[11]_net_1 ), .B(\cnt[13]_net_1 ), 
        .Y(state_tr0_0_a3_1));
    NOR3C \cnt_RNIU2GC2[4]  (.A(vd_stp_en_i_a3_4), .B(vd_stp_en_i_a3_3)
        , .C(N_73), .Y(vd_stp_en_i_a3_9));
    NOR3A \state_RNO_1[0]  (.A(state_tr0_0_a3_2), .B(\cnt[0]_net_1 ), 
        .C(\cnt[1]_net_1 ), .Y(state_tr0_0_a3_7));
    DFN1C0 \cnt[4]  (.D(N_20), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[4]_net_1 ));
    DFN1C0 \cnt[9]  (.D(cnt_n9), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[9]_net_1 ));
    NOR2A \cnt_RNO[0]  (.A(cs_i_1), .B(\cnt[0]_net_1 ), .Y(cnt_n0));
    OR3C \cnt_RNO_0[14]  (.A(\cnt[12]_net_1 ), .B(\cnt[13]_net_1 ), .C(
        cnt_N_13_mux), .Y(N_74));
    DFN1C0 \cnt[0]  (.D(cnt_n0), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[0]_net_1 ));
    NOR2B \cnt_RNI34RL_0[1]  (.A(\cnt[1]_net_1 ), .B(\cnt[0]_net_1 ), 
        .Y(cnt_m2_0_a2_0));
    NOR3B \cnt_RNO[4]  (.A(N_33), .B(cs_i_1), .C(N_97), .Y(N_20));
    NOR2 \state_RNO_4[0]  (.A(\cnt[10]_net_1 ), .B(\cnt[8]_net_1 ), .Y(
        state_tr0_0_a3_2));
    DFN1C0 \state[0]  (.D(\state_RNO_0[0]_net_1 ), .CLK(cur_clk), .CLR(
        n_rst_c), .Q(cs_i_1));
    XA1 \cnt_RNO[6]  (.A(cnt_N_7_mux_0_0), .B(\cnt[6]_net_1 ), .C(
        cs_i_1), .Y(\cnt_RNO_2[6]_net_1 ));
    NOR2B \cnt_RNI5JTG[11]  (.A(\cnt[11]_net_1 ), .B(\cnt[10]_net_1 ), 
        .Y(cnt_m6_0_a2_0));
    NOR2B \cnt_RNIBCRL[5]  (.A(\cnt[4]_net_1 ), .B(\cnt[5]_net_1 ), .Y(
        cnt_m5_0_a2_2));
    XA1 \cnt_RNO[15]  (.A(\cnt[15]_net_1 ), .B(cnt_N_3_mux_0), .C(
        cs_i_1), .Y(cnt_n15));
    XA1A \cnt_RNO[9]  (.A(\cnt[9]_net_1 ), .B(N_38), .C(cs_i_1), .Y(
        cnt_n9));
    GND GND_i (.Y(GND));
    NOR2B \cnt_RNO_5[10]  (.A(\cnt[8]_net_1 ), .B(\cnt[9]_net_1 ), .Y(
        cnt_m7_0_a2_1));
    NOR2 \cnt_RNI6KTG[10]  (.A(\cnt[10]_net_1 ), .B(\cnt[12]_net_1 ), 
        .Y(vd_stp_en_i_a3_2));
    DFN1C0 \cnt[13]  (.D(cnt_n13), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[13]_net_1 ));
    NOR3A \state_RNO_5[0]  (.A(state_tr0_0_a3_1), .B(\cnt[14]_net_1 ), 
        .C(\cnt[15]_net_1 ), .Y(state_tr0_0_a3_6));
    OR2A \cnt_RNO_0[9]  (.A(\cnt[8]_net_1 ), .B(N_36), .Y(N_38));
    OR3B \cnt_RNIV1KM1[4]  (.A(\cnt[3]_net_1 ), .B(\cnt[4]_net_1 ), .C(
        N_31), .Y(N_33));
    DFN1C0 \cnt[7]  (.D(N_14), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[7]_net_1 ));
    NOR3C \state_RNO_2[0]  (.A(state_tr0_0_a3_6), .B(cs_i_1), .C(
        state_tr0_0_a3_9), .Y(state_tr0_0_a3_12));
    OR2A \cnt_RNIMNO01[2]  (.A(\cnt[2]_net_1 ), .B(N_30), .Y(N_31));
    DFN1C0 \cnt[10]  (.D(cnt_n10), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[10]_net_1 ));
    NOR3C \cnt_RNO_1[11]  (.A(cnt_m6_0_a2_5_0), .B(\cnt[3]_net_1 ), .C(
        cnt_m5_0_a2_2), .Y(cnt_m6_0_a2_5_6));
    XA1A \cnt_RNO[5]  (.A(\cnt[5]_net_1 ), .B(N_33), .C(cs_i_1), .Y(
        N_18));
    DFN1C0 \cnt[3]  (.D(N_22), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[3]_net_1 ));
    NOR2B \cnt_RNO_2[11]  (.A(\cnt[10]_net_1 ), .B(\cnt[2]_net_1 ), .Y(
        cnt_m6_0_a2_5_0));
    NOR3 \cnt_RNI3IRR[15]  (.A(\cnt[14]_net_1 ), .B(\cnt[15]_net_1 ), 
        .C(\cnt[5]_net_1 ), .Y(vd_stp_en_i_a3_5));
    XA1A \cnt_RNO[14]  (.A(\cnt[14]_net_1 ), .B(N_74), .C(cs_i_1), .Y(
        cnt_n14));
    XNOR2 \cnt_RNO_1[10]  (.A(\cnt[10]_net_1 ), .B(\cnt[4]_net_1 ), .Y(
        \cnt_RNO_1[10]_net_1 ));
    NOR3C \cnt_RNO_4[10]  (.A(\cnt[7]_net_1 ), .B(\cnt[6]_net_1 ), .C(
        cnt_m7_0_a2_1), .Y(cnt_m7_0_a2_3));
    NOR3B \cnt_RNO_0[11]  (.A(cnt_m6_0_a2_5), .B(cnt_m6_0_a2_5_6), .C(
        N_30), .Y(cnt_N_13_mux_0));
    XA1 \cnt_RNO[11]  (.A(\cnt[11]_net_1 ), .B(cnt_N_13_mux_0), .C(
        cs_i_1), .Y(cnt_n11));
    OR2A \cnt_RNISTO01[4]  (.A(\cnt[4]_net_1 ), .B(N_103), .Y(N_73));
    NOR3B \cnt_RNO_2[10]  (.A(cnt_m7_0_a2_4), .B(cnt_m7_0_a2_3), .C(
        N_31), .Y(cnt_N_15_mux));
    OR3C \state_RNO[0]  (.A(state_tr0_0_a3_8), .B(state_tr0_0_a3_7), 
        .C(state_tr0_0_a3_12), .Y(\state_RNO_0[0]_net_1 ));
    MX2B \cnt_RNO[10]  (.A(d_N_3_mux_3), .B(\cnt_RNO_1[10]_net_1 ), .S(
        cnt_N_15_mux), .Y(cnt_n10));
    DFN1C0 \cnt[15]  (.D(cnt_n15), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[15]_net_1 ));
    NOR2B \cnt_RNO_1[6]  (.A(\cnt[2]_net_1 ), .B(\cnt[5]_net_1 ), .Y(
        cnt_m2_0_a2_1));
    OR2B \cnt_RNI34RL[1]  (.A(\cnt[1]_net_1 ), .B(\cnt[0]_net_1 ), .Y(
        N_30));
    AO1B \state_RNIST2M4[0]  (.A(vd_stp_en_i_a3_9), .B(
        vd_stp_en_i_a3_8), .C(cs_i_1), .Y(N_29));
    NOR2B \cnt_RNO_0[10]  (.A(\cnt[10]_net_1 ), .B(cs_i_1), .Y(
        d_N_3_mux_3));
    NOR3C \cnt_RNICGFC2[2]  (.A(cnt_m5_0_a2_2), .B(cnt_m5_0_a2_1), .C(
        cnt_m5_0_a2_3), .Y(cnt_N_11_mux_2));
    NOR2 \state_RNO_3[0]  (.A(\cnt[9]_net_1 ), .B(\cnt[12]_net_1 ), .Y(
        state_tr0_0_a3_4));
    DFN1C0 \cnt[5]  (.D(N_18), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[5]_net_1 ));
    INV \state_RNIDURB[0]  (.A(cs_i_1), .Y(cs_i_1_i));
    XA1A \cnt_RNO[13]  (.A(\cnt[13]_net_1 ), .B(N_72), .C(cs_i_1), .Y(
        cnt_n13));
    NOR3C \cnt_RNI4KMH1[3]  (.A(cnt_m6_0_a2_0), .B(\cnt[3]_net_1 ), .C(
        cnt_m5_0_a2_2), .Y(cnt_m6_0_a2_6));
    XA1 \cnt_RNO[12]  (.A(\cnt[12]_net_1 ), .B(cnt_N_13_mux), .C(
        cs_i_1), .Y(cnt_n12));
    DFN1C0 \cnt[12]  (.D(cnt_n12), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[12]_net_1 ));
    XA1 \cnt_RNO[7]  (.A(\cnt[7]_net_1 ), .B(cnt_N_11_mux_2), .C(
        cs_i_1), .Y(N_14));
    DFN1C0 \cnt[14]  (.D(cnt_n14), .CLK(cur_clk), .CLR(n_rst_c), .Q(
        \cnt[14]_net_1 ));
    NOR2B \cnt_RNINOO01[3]  (.A(\cnt[3]_net_1 ), .B(cnt_m2_0_a2_0), .Y(
        cnt_m5_0_a2_3));
    
endmodule


module spi_rx_12s_0(
       cur_vd,
       vd_done,
       cs_i_1_i,
       cur_clk,
       n_rst_c,
       din_12_c
    );
output [11:0] cur_vd;
output vd_done;
output cs_i_1_i;
input  cur_clk;
input  n_rst_c;
input  din_12_c;

    wire N_29, cs_i_1, GND, VCC;
    
    spi_stp_12s_1_1 VD_STP (.cur_vd({cur_vd[11], cur_vd[10], cur_vd[9], 
        cur_vd[8], cur_vd[7], cur_vd[6], cur_vd[5], cur_vd[4], 
        cur_vd[3], cur_vd[2], cur_vd[1], cur_vd[0]}), .N_29(N_29), 
        .din_12_c(din_12_c), .n_rst_c(n_rst_c), .cur_clk(cur_clk));
    sig_gen_10_0 SPI_RDYSIG (.cs_i_1(cs_i_1), .n_rst_c(n_rst_c), 
        .cur_clk(cur_clk), .vd_done(vd_done));
    VCC VCC_i (.Y(VCC));
    spi_ctl_12s_0 SPICTL (.n_rst_c(n_rst_c), .cur_clk(cur_clk), .N_29(
        N_29), .cs_i_1(cs_i_1), .cs_i_1_i(cs_i_1_i));
    GND GND_i (.Y(GND));
    
endmodule


module integral_calc_13s_0_4(
       sr_new,
       sr_old,
       sr_new_1_0,
       sr_new_0_0,
       integral,
       integral_i,
       integral_0_0,
       integral_1_0,
       calc_int,
       N_46_1,
       n_rst_c,
       clk_c
    );
input  [12:0] sr_new;
input  [12:0] sr_old;
input  sr_new_1_0;
input  sr_new_0_0;
output [25:6] integral;
output [25:24] integral_i;
output integral_0_0;
output integral_1_0;
input  calc_int;
output N_46_1;
input  n_rst_c;
input  clk_c;

    wire \un1_integ[25] , \un1_next_int_0_iv_0[13] , next_int_1_sqmuxa, 
        next_int_0_sqmuxa_1, N_46_1_0, \state[0]_net_1 , 
        \state[1]_net_1 , N_12, N_10, \DWACT_FINC_E[0] , N_5, 
        \DWACT_FINC_E[4] , N_2, \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , 
        N_12_0, N_10_0, \DWACT_FINC_E_0[0] , N_5_0, 
        \DWACT_FINC_E_0[4] , N_2_0, \DWACT_FINC_E_0[7] , 
        \DWACT_FINC_E_0[6] , ADD_26x26_fast_I255_Y_0, 
        \un1_next_int_0_iv[13] , ADD_26x26_fast_I254_Y_0, 
        ADD_26x26_fast_I253_Y_0, ADD_26x26_fast_I252_Y_0, 
        ADD_26x26_fast_I247_Y_0, ADD_26x26_fast_I204_Y_3, N502, N517, 
        ADD_26x26_fast_I204_Y_2, N398, ADD_26x26_fast_I204_Y_0, N455, 
        ADD_26x26_fast_I205_Y_3, N504, N519, ADD_26x26_fast_I205_Y_2, 
        N457, N450, ADD_26x26_fast_I205_Y_1, ADD_26x26_fast_I205_Y_0, 
        N400, ADD_26x26_fast_I250_Y_0, ADD_26x26_fast_I251_Y_0, 
        ADD_26x26_fast_I206_Y_2, ADD_26x26_fast_I206_un1_Y_0, N522, 
        ADD_26x26_fast_I206_Y_1, N402, N459, ADD_26x26_fast_I245_Y_0, 
        ADD_26x26_fast_I207_Y_2, ADD_26x26_fast_I207_un1_Y_0, N524, 
        ADD_26x26_fast_I207_Y_1, N461, N454, ADD_26x26_fast_I207_Y_0, 
        N404, ADD_26x26_fast_I210_Y_0, N467, N460, 
        ADD_26x26_fast_I212_Y_0, N533, N518, ADD_26x26_fast_I244_Y_0, 
        ADD_26x26_fast_I243_Y_0, ADD_26x26_fast_I242_Y_0, 
        \un1_next_int[12] , ADD_26x26_fast_I208_Y_1, 
        ADD_26x26_fast_I208_un1_Y_0, N526, ADD_26x26_fast_I208_Y_0, 
        N463, N456, ADD_26x26_fast_I209_Y_1, 
        ADD_26x26_fast_I209_un1_Y_0, N528, ADD_26x26_fast_I209_Y_0, 
        N465, N458, ADD_26x26_fast_I211_Y_0, N469, N462, 
        ADD_26x26_fast_I204_un1_Y_0, ADD_26x26_fast_I239_Y_0, 
        \un2_next_int_m[9] , \un1_next_int_iv_1[9] , 
        ADD_26x26_fast_I212_un1_Y_0, N480, N488, N442, 
        ADD_26x26_fast_I213_un1_Y_0, N482, N490, \un1_next_int[0] , 
        ADD_26x26_fast_I211_Y_1_0, N470, N506, N537, N543, N512, N487, 
        I162_un1_Y, N510, N485, I161_un1_Y, N508, 
        ADD_26x26_fast_I237_Y_0, \un2_next_int_m[7] , 
        \un1_next_int_iv_1[7] , ADD_26x26_fast_I236_Y_0, 
        \un1_next_int[6] , ADD_26x26_fast_I235_Y_0, 
        \un2_next_int_m[5] , \un1_next_int_iv_1[5] , \integ[5]_net_1 , 
        ADD_26x26_fast_I232_Y_0, \integ[2]_net_1 , \un1_next_int[2] , 
        ADD_26x26_fast_I125_Y_0, ADD_26x26_fast_I79_Y_0, 
        \un1_next_int_iv_0[10] , \inf_abs1[10]_net_1 , 
        \un1_next_int_iv_0[11] , \inf_abs1[11]_net_1 , 
        \un1_next_int_iv_0[7] , \inf_abs0_m[7] , \inf_abs1[7]_net_1 , 
        \un1_next_int_iv_0[8] , \inf_abs1[8]_net_1 , 
        \un1_next_int_iv_1[6] , \un1_next_int_iv_0[6] , 
        \inf_abs0_m[6] , \inf_abs1[6]_net_1 , \inf_abs0_m[9] , 
        \un18_next_int_m[9] , \inf_abs1_m[9] , \un1_next_int_iv_0[12] , 
        \inf_abs1_a_1[12] , \un1_next_int_iv_0[0] , 
        \inf_abs1[0]_net_1 , \inf_abs0_m[5] , \un18_next_int_m[5] , 
        \inf_abs1_m[5] , \un1_next_int_iv_1[4] , \inf_abs1_m[4] , 
        \un1_next_int_iv_0[4] , \un18_next_int_m[4] , \inf_abs0_m[4] , 
        \un1_next_int_iv_1[3] , \inf_abs1_m[3] , \un18_next_int_m[3] , 
        \inf_abs0_m[3] , \un1_next_int_iv_0[2] , \inf_abs1[2]_net_1 , 
        \un1_next_int_iv_1[1] , \un18_next_int_m[1] , \inf_abs1_m[1] , 
        \un2_next_int_m[1] , \un1_next_int[3] , \un2_next_int_m[3] , 
        \un1_integ[5] , \un1_integ[9] , I194_un1_Y, \un1_integ[21] , 
        I176_un1_Y, \un1_integ[15] , N521, I188_un1_Y, \un1_integ[13] , 
        N525, I190_un1_Y, \un1_integ[3] , \integ[3]_net_1 , N491, 
        \un1_next_int[1] , \inf_abs0_m[1] , \un2_next_int_m[12] , N399, 
        I204_un1_Y, \un1_next_int[11] , \inf_abs0_m[11] , 
        \un2_next_int_m[11] , \un1_integ[11] , N649, \un1_integ[7] , 
        I212_un1_Y, N403, \un1_integ[23] , I172_un1_Y, \un1_integ[0] , 
        N_3, \integ[0]_net_1 , \un1_integ[17] , N401, 
        \un1_next_int[4] , \un2_next_int_m[4] , \un1_integ[1] , 
        \integ[1]_net_1 , \un1_integ[4] , \integ[4]_net_1 , I205_un1_Y, 
        N520, N658, N631, ADD_26x26_fast_I211_Y_1_tz, \un1_integ[22] , 
        I174_un1_Y, \un1_integ[18] , \un1_integ[24] , \un1_integ[12] , 
        N527, I191_un1_Y, \un1_integ[6] , \un1_integ[14] , N523, 
        I189_un1_Y, \un1_integ[16] , N635, \un1_integ[19] , N629, 
        \un1_integ[2] , N493, \un1_integ[10] , \un1_next_int[10] , 
        N652, \un1_integ[20] , I178_un1_Y, \un1_integ[8] , 
        \un1_next_int[8] , \inf_abs0_m[0] , \un2_next_int_m[0] , 
        \inf_abs0_m[2] , \un2_next_int_m[2] , \un2_next_int_m[6] , 
        \inf_abs0_m[8] , \un2_next_int_m[8] , \inf_abs0_m[10] , 
        \un2_next_int_m[10] , I180_un1_Y, I210_un1_Y, N514, N530, 
        I186_un1_Y, I213_un1_Y, N477, I154_un1_Y, 
        ADD_26x26_fast_I211_un1_Y_0, N478, N486, N474, I158_un1_Y, 
        N489, I163_un1_Y, N481, I195_un1_Y, N431, N333, N336, N473, 
        N424, N421, N420, N425, N345, N342, I146_un1_Y, N417, N416, 
        N339, N466, I118_un1_Y, N436, N440, N437, N441, I110_un1_Y, 
        N428, N335, N338, N432, N430, N332, N468, N475, I152_un1_Y, 
        N433, N347, N348, I114_un1_Y, I121_un1_Y, I193_un1_Y, N341, 
        \inf_abs0[6]_net_1 , \inf_abs0[7]_net_1 , \inf_abs0[8]_net_1 , 
        \inf_abs0[10]_net_1 , \state_RNO_0[1] , \inf_abs0_a_0[6] , 
        \inf_abs0_a_0[7] , \inf_abs0_a_0[8] , \inf_abs0_a_0[10] , 
        \inf_abs1_a_1[6] , \inf_abs1_a_1[7] , \inf_abs1_a_1[8] , 
        \inf_abs1_a_1[10] , \inf_abs0[0]_net_1 , \inf_abs0[2]_net_1 , 
        \inf_abs0_a_0[2] , \inf_abs1_a_1[2] , \state_RNO[0]_net_1 , 
        N413, I150_un1_Y, \inf_abs1_a_1[4] , \inf_abs0_a_0[4] , N329, 
        N321, N320, N405, N406, N412, N410, N409, N408, N317, N357, 
        N354, N414, N418, N415, N318, N407, N464, N411, N353, 
        \inf_abs1_a_1[11] , \inf_abs0[11]_net_1 , \inf_abs0_a_0[11] , 
        N351, N350, I192_un1_Y, N484, N483, N476, N435, N327, N434, 
        N326, \inf_abs0_a_0[9] , \inf_abs1_a_1[9] , \inf_abs0_a_0[12] , 
        \inf_abs0_a_0[1] , \inf_abs1_a_1[1] , N344, \inf_abs1_a_1[5] , 
        \inf_abs0_a_0[5] , \inf_abs1_a_1[3] , \inf_abs0_a_0[3] , N422, 
        N438, N472, I148_un1_Y, N471, N479, N439, N423, N419, 
        I68_un1_Y, I108_un1_Y, N426, N_3_0, \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[5] , N_4, \DWACT_FINC_E[3] , N_6, N_7, N_8, 
        \DWACT_FINC_E[1] , N_9, N_11, N_3_1, \DWACT_FINC_E_0[2] , 
        \DWACT_FINC_E_0[5] , N_4_0, \DWACT_FINC_E_0[3] , N_6_0, N_7_0, 
        N_8_0, \DWACT_FINC_E_0[1] , N_9_0, N_11_0, GND, VCC;
    
    AO1 un1_integ_0_0_ADD_26x26_fast_I56_Y (.A(N341), .B(N345), .C(
        N344), .Y(N424));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I148_un1_Y (.A(N479), .B(N472), 
        .Y(I148_un1_Y));
    NOR2 inf_abs1_a_1_I_15 (.A(sr_old[3]), .B(sr_old[4]), .Y(
        \DWACT_FINC_E[1] ));
    XNOR2 inf_abs1_a_1_I_23 (.A(sr_old[8]), .B(N_6), .Y(
        \inf_abs1_a_1[8] ));
    DFN1C0 \state[0]  (.D(\state_RNO[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[0]_net_1 ));
    XNOR2 inf_abs1_a_1_I_17 (.A(sr_old[6]), .B(N_8), .Y(
        \inf_abs1_a_1[6] ));
    DFN1E0C0 \integ[13]  (.D(\un1_integ[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[13]));
    DFN1E0C0 \integ[24]  (.D(\un1_integ[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[24]));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I245_Y_0 (.A(integral[15]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I245_Y_0));
    NOR2A \state_RNIRATB[0]  (.A(\state[0]_net_1 ), .B(sr_new[12]), .Y(
        next_int_1_sqmuxa));
    OR3 un1_integ_0_0_ADD_26x26_fast_I7_P0N (.A(\un2_next_int_m[7] ), 
        .B(\un1_next_int_iv_1[7] ), .C(integral[7]), .Y(N339));
    NOR3B inf_abs0_a_0_I_19 (.A(\DWACT_FINC_E_0[2] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[6]), .Y(N_7_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I172_un1_Y (.A(N506), .B(N521), 
        .Y(I172_un1_Y));
    NOR3B inf_abs0_a_0_I_16 (.A(\DWACT_FINC_E_0[1] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[5]), .Y(N_8_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I41_Y (.A(integral[16]), .B(
        integral[17]), .C(\un1_next_int_0_iv_0[13] ), .Y(N409));
    OA1 un1_integ_0_0_ADD_26x26_fast_I204_un1_Y (.A(N533), .B(
        I194_un1_Y), .C(ADD_26x26_fast_I204_un1_Y_0), .Y(I204_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I86_Y (.A(N408), .B(N404), .Y(
        N457));
    AO1 un1_integ_0_0_ADD_26x26_fast_I98_Y (.A(N420), .B(N417), .C(
        N416), .Y(N469));
    INV \integ_RNIFIQB[25]  (.A(integral[25]), .Y(integral_i[25]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I176_un1_Y (.A(N510), .B(N525), 
        .Y(I176_un1_Y));
    OR3 un1_integ_0_0_ADD_26x26_fast_I193_Y (.A(N477), .B(I154_un1_Y), 
        .C(I193_un1_Y), .Y(N652));
    NOR3B \state_RNIRDV13[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[8]_net_1 ), .Y(\un2_next_int_m[8] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I158_un1_Y (.A(N489), .B(N482), 
        .Y(I158_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I150_un1_Y (.A(N481), .B(N474), 
        .Y(I150_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I51_Y (.A(N354), .B(N351), .Y(
        N419));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I230_Y (.A(N_3), .B(
        \integ[0]_net_1 ), .C(\un1_next_int[0] ), .Y(\un1_integ[0] ));
    NOR3A \state_RNITH3C[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), .C(
        sr_old[9]), .Y(\un18_next_int_m[9] ));
    OR2 \state_RNIQ6VM2[0]  (.A(\un1_next_int_iv_1[3] ), .B(
        \un2_next_int_m[3] ), .Y(\un1_next_int[3] ));
    NOR2B inf_abs1_a_1_I_34 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .Y(N_2_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I253_Y (.A(I172_un1_Y), .B(
        ADD_26x26_fast_I206_Y_2), .C(ADD_26x26_fast_I253_Y_0), .Y(
        \un1_integ[23] ));
    DFN1E0C0 \integ[21]  (.D(\un1_integ[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[21]));
    XNOR2 inf_abs1_a_1_I_7 (.A(sr_old[2]), .B(N_12_0), .Y(
        \inf_abs1_a_1[2] ));
    DFN1E0C0 \integ_1[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral_1_0));
    OR2 \state_RNIGQRN[1]  (.A(next_int_1_sqmuxa), .B(
        next_int_0_sqmuxa_1), .Y(\un1_next_int_0_iv_0[13] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I190_un1_Y (.A(N487), .B(
        I162_un1_Y), .C(N526), .Y(I190_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I146_Y (.A(I146_un1_Y), .B(N469), 
        .Y(N523));
    AO1 un1_integ_0_0_ADD_26x26_fast_I142_Y (.A(N473), .B(N466), .C(
        N465), .Y(N519));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I244_Y_0 (.A(integral[14]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I244_Y_0));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I231_Y (.A(\un1_next_int[1] ), 
        .B(\integ[1]_net_1 ), .C(N442), .Y(\un1_integ[1] ));
    OR2 \state_RNI9OIT2[0]  (.A(\un1_next_int_iv_1[4] ), .B(
        \un2_next_int_m[4] ), .Y(\un1_next_int[4] ));
    AND3 inf_abs1_a_1_I_24 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E_0[4] ));
    XNOR2 inf_abs1_a_1_I_32 (.A(sr_old[11]), .B(N_3_0), .Y(
        \inf_abs1_a_1[11] ));
    DFN1E0C0 \integ[15]  (.D(\un1_integ[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[15]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I213_un1_Y (.A(
        ADD_26x26_fast_I213_un1_Y_0), .B(N520), .Y(I213_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I103_Y (.A(N421), .B(N425), .Y(
        N474));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I125_Y (.A(N399), .B(
        ADD_26x26_fast_I125_Y_0), .C(N456), .Y(N502));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_1 (.A(
        ADD_26x26_fast_I209_un1_Y_0), .B(N528), .C(
        ADD_26x26_fast_I209_Y_0), .Y(ADD_26x26_fast_I209_Y_1));
    OR3 \state_RNI0GCN1[0]  (.A(\un18_next_int_m[1] ), .B(
        \inf_abs1_m[1] ), .C(\un2_next_int_m[1] ), .Y(
        \un1_next_int_iv_1[1] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I97_Y (.A(N415), .B(N419), .Y(
        N468));
    AO1 un1_integ_0_0_ADD_26x26_fast_I94_Y (.A(N416), .B(N413), .C(
        N412), .Y(N465));
    NOR2 inf_abs0_a_0_I_6 (.A(sr_new[0]), .B(sr_new[1]), .Y(N_12));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I151_Y (.A(N482), .B(N474), .Y(
        N528));
    AND3 inf_abs1_a_1_I_22 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_6));
    AO1 un1_integ_0_0_ADD_26x26_fast_I74_Y (.A(N318), .B(
        \un1_next_int[0] ), .C(N317), .Y(N442));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I238_Y (.A(\un1_next_int[8] ), 
        .B(integral[8]), .C(N658), .Y(\un1_integ[8] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I121_Y (.A(I121_un1_Y), .B(N440), 
        .Y(N493));
    NOR3 inf_abs0_a_0_I_10 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2])
        , .Y(\DWACT_FINC_E[0] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I154_un1_Y (.A(N485), .B(N478), 
        .Y(I154_un1_Y));
    OR3 un1_integ_0_0_ADD_26x26_fast_I5_P0N (.A(\un2_next_int_m[5] ), 
        .B(\un1_next_int_iv_1[5] ), .C(\integ[5]_net_1 ), .Y(N333));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I236_Y_0 (.A(integral[6]), .B(
        \un1_next_int[6] ), .Y(ADD_26x26_fast_I236_Y_0));
    XA1A \state_RNISL511[1]  (.A(sr_old[12]), .B(\inf_abs1[11]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[11] ));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I246_Y (.A(
        \un1_next_int_0_iv_0[13] ), .B(integral[16]), .C(N635), .Y(
        \un1_integ[16] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I252_Y_0 (.A(integral[22]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I252_Y_0));
    MX2 \inf_abs0[6]  (.A(sr_new[6]), .B(\inf_abs0_a_0[6] ), .S(
        sr_new_1_0), .Y(\inf_abs0[6]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I39_Y (.A(integral[18]), .B(
        integral[17]), .C(\un1_next_int_0_iv[13] ), .Y(N407));
    OA1B un1_integ_0_0_ADD_26x26_fast_I32_Y (.A(integral[20]), .B(
        integral[21]), .C(\un1_next_int_0_iv_0[13] ), .Y(N400));
    OR3 un1_integ_0_0_ADD_26x26_fast_I213_Y (.A(I186_un1_Y), .B(N519), 
        .C(I213_un1_Y), .Y(N635));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I194_un1_Y (.A(N480), .B(N488), 
        .C(N442), .Y(I194_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I108_un1_Y (.A(N339), .B(N342), 
        .C(N430), .Y(I108_un1_Y));
    NOR2A inf_abs0_a_0_I_11 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .Y(
        N_10));
    AO1B un1_integ_0_0_ADD_26x26_fast_I125_Y_0 (.A(integral[23]), .B(
        integral[24]), .C(\un1_next_int_0_iv_0[13] ), .Y(
        ADD_26x26_fast_I125_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I211_Y_1_0 (.A(N462), .B(N470), 
        .Y(ADD_26x26_fast_I211_Y_1_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I100_Y (.A(N422), .B(N419), .C(
        N418), .Y(N471));
    OR2 un1_integ_0_0_ADD_26x26_fast_I12_P0N (.A(\un1_next_int[12] ), 
        .B(integral[12]), .Y(N354));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I10_G0N (.A(\un1_next_int[10] ), 
        .B(integral[10]), .Y(N347));
    OR2 \state_RNI2AO92[0]  (.A(\un1_next_int_iv_1[1] ), .B(
        \inf_abs0_m[1] ), .Y(\un1_next_int[1] ));
    DFN1E0C0 \integ[12]  (.D(\un1_integ[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[12]));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I109_Y (.A(N339), .B(N342), .C(
        N431), .Y(N480));
    XNOR2 inf_abs1_a_1_I_35 (.A(sr_old[12]), .B(N_2_0), .Y(
        \inf_abs1_a_1[12] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I205_Y_0 (.A(integral[22]), .B(
        integral[23]), .C(\un1_next_int_0_iv_0[13] ), .Y(
        ADD_26x26_fast_I205_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I115_Y (.A(N437), .B(N433), .Y(
        N486));
    NOR2B \state_RNIUKRC[1]  (.A(\inf_abs1_a_1[5] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[5] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I12_G0N (.A(\un1_next_int[12] ), 
        .B(integral[12]), .Y(N353));
    OR3 \state_RNII11B1[1]  (.A(\inf_abs1_m[3] ), .B(
        \un18_next_int_m[3] ), .C(\inf_abs0_m[3] ), .Y(
        \un1_next_int_iv_1[3] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_0 (.A(N463), .B(N456), .C(
        N455), .Y(ADD_26x26_fast_I208_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I111_Y (.A(N339), .B(N336), .C(
        N433), .Y(N482));
    NOR2A inf_abs1_a_1_I_25 (.A(\DWACT_FINC_E_0[4] ), .B(sr_old[8]), 
        .Y(N_5_0));
    OR3 \state_RNIJS7S7[0]  (.A(\inf_abs0_m[11] ), .B(
        \un1_next_int_iv_0[11] ), .C(\un2_next_int_m[11] ), .Y(
        \un1_next_int[11] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I250_Y_0 (.A(integral[20]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I250_Y_0));
    NOR3A inf_abs1_a_1_I_27 (.A(\DWACT_FINC_E_0[4] ), .B(sr_old[8]), 
        .C(sr_old[9]), .Y(N_4));
    DFN1E0C0 \integ[10]  (.D(\un1_integ[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[10]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I188_un1_Y (.A(N522), .B(N537), 
        .Y(I188_un1_Y));
    OA1 un1_integ_0_0_ADD_26x26_fast_I180_un1_Y (.A(N475), .B(
        I152_un1_Y), .C(N514), .Y(I180_un1_Y));
    XA1A \state_RNI89FH[1]  (.A(sr_old[12]), .B(\inf_abs1[2]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[2] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I6_G0N (.A(\un1_next_int[6] ), 
        .B(integral[6]), .Y(N335));
    MX2 \inf_abs1[10]  (.A(sr_old[10]), .B(\inf_abs1_a_1[10] ), .S(
        sr_old[12]), .Y(\inf_abs1[10]_net_1 ));
    NOR2B \state_RNINPHC[1]  (.A(\inf_abs1_a_1[3] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[3] ));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I249_Y (.A(
        \un1_next_int_0_iv_0[13] ), .B(integral[19]), .C(N629), .Y(
        \un1_integ[19] ));
    GND GND_i (.Y(GND));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I146_un1_Y (.A(N477), .B(N470), 
        .Y(I146_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I6_P0N (.A(\un1_next_int[6] ), .B(
        integral[6]), .Y(N336));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I68_un1_Y (.A(\integ[2]_net_1 ), 
        .B(\un1_next_int[2] ), .C(N327), .Y(I68_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I212_un1_Y_0 (.A(N480), .B(N488)
        , .C(N442), .Y(ADD_26x26_fast_I212_un1_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I1_G0N (.A(\un1_next_int[1] ), 
        .B(\integ[1]_net_1 ), .Y(N320));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I107_Y (.A(N339), .B(N336), .C(
        N425), .Y(N478));
    XNOR2 inf_abs1_a_1_I_9 (.A(sr_old[3]), .B(N_11), .Y(
        \inf_abs1_a_1[3] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I38_Y (.A(integral[17]), .B(
        integral[18]), .C(\un1_next_int_0_iv[13] ), .Y(N406));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I209_un1_Y_0 (.A(N543), .B(N512)
        , .Y(ADD_26x26_fast_I209_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_3 (.A(N504), .B(N519), .C(
        ADD_26x26_fast_I205_Y_2), .Y(ADD_26x26_fast_I205_Y_3));
    AX1D un1_integ_0_0_ADD_26x26_fast_I255_Y (.A(I204_un1_Y), .B(
        ADD_26x26_fast_I204_Y_3), .C(ADD_26x26_fast_I255_Y_0), .Y(
        \un1_integ[25] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I204_Y_0 (.A(integral[24]), .B(
        integral[23]), .C(\un1_next_int_0_iv_0[13] ), .Y(
        ADD_26x26_fast_I204_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I243_Y (.A(N525), .B(I190_un1_Y), 
        .C(ADD_26x26_fast_I243_Y_0), .Y(\un1_integ[13] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I69_Y (.A(\integ[2]_net_1 ), .B(
        \un1_next_int[2] ), .C(N327), .Y(N437));
    AO1 un1_integ_0_0_ADD_26x26_fast_I62_Y (.A(N332), .B(N336), .C(
        N335), .Y(N430));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I193_un1_Y (.A(N478), .B(N486), 
        .C(N493), .Y(I193_un1_Y));
    NOR3B \state_RNIA4OB3[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[10]_net_1 ), .Y(\un2_next_int_m[10] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I153_Y (.A(N484), .B(N476), .Y(
        N530));
    NOR2B \state_RNILFUB[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), .Y(
        next_int_0_sqmuxa_1));
    NOR3B \state_RNIS9H53[0]  (.A(sr_new_1_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[12] ), .Y(\un2_next_int_m[12] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I152_un1_Y (.A(N483), .B(N476), 
        .Y(I152_un1_Y));
    OA1A \state_RNIB68S[1]  (.A(sr_old[12]), .B(\inf_abs1_a_1[12] ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[12] ));
    XNOR2 inf_abs0_a_0_I_7 (.A(sr_new[2]), .B(N_12), .Y(
        \inf_abs0_a_0[2] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I7_G0N (.A(\un2_next_int_m[7] ), 
        .B(\un1_next_int_iv_1[7] ), .C(integral[7]), .Y(N338));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I49_Y (.A(N357), .B(N354), .Y(
        N417));
    OA1B un1_integ_0_0_ADD_26x26_fast_I42_Y (.A(integral[16]), .B(
        integral[15]), .C(\un1_next_int_0_iv_0[13] ), .Y(N410));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I145_Y (.A(N468), .B(N476), .Y(
        N522));
    XA1A \state_RNI97DI[1]  (.A(sr_old[12]), .B(\inf_abs1[8]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[8] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I10_P0N (.A(\un1_next_int[10] ), 
        .B(integral[10]), .Y(N348));
    OR2 un1_integ_0_0_ADD_26x26_fast_I1_P0N (.A(\un1_next_int[1] ), .B(
        \integ[1]_net_1 ), .Y(N321));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I192_un1_Y (.A(N530), .B(N491), 
        .Y(I192_un1_Y));
    NOR3A \state_RNIPD3C[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), .C(
        sr_old[5]), .Y(\un18_next_int_m[5] ));
    NOR3A inf_abs0_a_0_I_13 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .C(
        sr_new[4]), .Y(N_9_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I141_Y (.A(N464), .B(N472), .Y(
        N518));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I93_Y (.A(N411), .B(N415), .Y(
        N464));
    AO1B un1_integ_0_0_ADD_26x26_fast_I37_Y (.A(integral[19]), .B(
        integral[18]), .C(\un1_next_int_0_iv[13] ), .Y(N405));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I0_G0N (.A(N_3), .B(
        \integ[0]_net_1 ), .Y(N317));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I73_Y (.A(N318), .B(N321), .Y(
        N441));
    AO1 un1_integ_0_0_ADD_26x26_fast_I52_Y (.A(N347), .B(N351), .C(
        N350), .Y(N420));
    NOR2A \state_RNO[1]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 ), 
        .Y(\state_RNO_0[1] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I34_Y (.A(integral[20]), .B(
        integral[19]), .C(\un1_next_int_0_iv[13] ), .Y(N402));
    AX1D un1_integ_0_0_ADD_26x26_fast_I236_Y (.A(N485), .B(I161_un1_Y), 
        .C(ADD_26x26_fast_I236_Y_0), .Y(\un1_integ[6] ));
    OR2 \state_RNIT9FU[1]  (.A(\un18_next_int_m[4] ), .B(
        \inf_abs0_m[4] ), .Y(\un1_next_int_iv_0[4] ));
    NOR3B \state_RNIN31V[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), .C(
        \inf_abs0_a_0[1] ), .Y(\un2_next_int_m[1] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I205_Y_1 (.A(
        ADD_26x26_fast_I205_Y_0), .B(N400), .Y(ADD_26x26_fast_I205_Y_1)
        );
    OR2 un1_integ_0_0_ADD_26x26_fast_I150_Y (.A(I150_un1_Y), .B(N473), 
        .Y(N527));
    XA1A \state_RNI158I[1]  (.A(sr_old[12]), .B(\inf_abs1[7]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[7] ));
    DFN1E0C0 \integ[0]  (.D(\un1_integ[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(\integ[0]_net_1 ));
    NOR2B \state_RNI2QBI[0]  (.A(sr_new[1]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[1] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I120_Y (.A(N439), .B(N442), .C(
        N438), .Y(N491));
    AO1 un1_integ_0_0_ADD_26x26_fast_I104_Y (.A(N423), .B(N426), .C(
        N422), .Y(N475));
    VCC VCC_i (.Y(VCC));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I129_Y (.A(N403), .B(N399), .C(
        N460), .Y(N506));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I113_Y (.A(N431), .B(N435), .Y(
        N484));
    MX2 \inf_abs0[0]  (.A(sr_new[0]), .B(sr_new[0]), .S(sr_new_1_0), 
        .Y(\inf_abs0[0]_net_1 ));
    OR2 \state_RNIN06B1[1]  (.A(\inf_abs1_m[4] ), .B(
        \un1_next_int_iv_0[4] ), .Y(\un1_next_int_iv_1[4] ));
    XNOR2 inf_abs0_a_0_I_28 (.A(sr_new[10]), .B(N_4_0), .Y(
        \inf_abs0_a_0[10] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I89_Y (.A(N411), .B(N407), .Y(
        N460));
    OR2 un1_integ_0_0_ADD_26x26_fast_I68_Y (.A(I68_un1_Y), .B(N326), 
        .Y(N436));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_0 (.A(N469), .B(N462), .C(
        N461), .Y(ADD_26x26_fast_I211_Y_0));
    DFN1E0C0 \integ[4]  (.D(\un1_integ[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(\integ[4]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I108_Y (.A(I108_un1_Y), .B(N426), 
        .Y(N479));
    NOR3 inf_abs1_a_1_I_18 (.A(sr_old[4]), .B(sr_old[3]), .C(sr_old[5])
        , .Y(\DWACT_FINC_E[2] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I3_G0N (.A(\un1_next_int[3] ), 
        .B(\integ[3]_net_1 ), .Y(N326));
    AO13 un1_integ_0_0_ADD_26x26_fast_I48_Y (.A(integral[13]), .B(N353)
        , .C(\un1_next_int_0_iv_0[13] ), .Y(N416));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I195_un1_Y (.A(N482), .B(N490), 
        .C(\un1_next_int[0] ), .Y(I195_un1_Y));
    DFN1E0C0 \integ[3]  (.D(\un1_integ[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(\integ[3]_net_1 ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I252_Y (.A(I174_un1_Y), .B(
        ADD_26x26_fast_I207_Y_2), .C(ADD_26x26_fast_I252_Y_0), .Y(
        \un1_integ[22] ));
    DFN1E0C0 \integ[6]  (.D(\un1_integ[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(integral[6]));
    XNOR2 inf_abs0_a_0_I_14 (.A(sr_new[5]), .B(N_9_0), .Y(
        \inf_abs0_a_0[5] ));
    AND3 inf_abs0_a_0_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[5] ), .Y(
        \DWACT_FINC_E[6] ));
    OR2 \state_RNI7GP14[0]  (.A(\un1_next_int_iv_0[12] ), .B(
        \un2_next_int_m[12] ), .Y(\un1_next_int[12] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y (.A(N533), .B(I194_un1_Y), 
        .C(ADD_26x26_fast_I239_Y_0), .Y(\un1_integ[9] ));
    NOR2 \state_RNI5T1E_0[0]  (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(N_46_1_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I58_Y (.A(N338), .B(N342), .C(
        N341), .Y(N426));
    OA1 un1_integ_0_0_ADD_26x26_fast_I67_Y (.A(\integ[4]_net_1 ), .B(
        \un1_next_int[4] ), .C(N327), .Y(N435));
    XNOR2 inf_abs0_a_0_I_12 (.A(sr_new[4]), .B(N_10), .Y(
        \inf_abs0_a_0[4] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I253_Y_0 (.A(integral[23]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I253_Y_0));
    OR3 \state_RNIKKJ73[0]  (.A(\inf_abs0_m[0] ), .B(
        \un1_next_int_iv_0[0] ), .C(\un2_next_int_m[0] ), .Y(
        \un1_next_int[0] ));
    NOR2B \state_RNIK28C[1]  (.A(\inf_abs1_a_1[1] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[1] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I64_Y (.A(N329), .B(N333), .C(
        N332), .Y(N432));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I204_un1_Y_0 (.A(N502), .B(N518)
        , .Y(ADD_26x26_fast_I204_un1_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I212_un1_Y (.A(
        ADD_26x26_fast_I212_un1_Y_0), .B(N518), .Y(I212_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I127_Y (.A(N450), .B(N458), .Y(
        N504));
    OR2 un1_integ_0_0_ADD_26x26_fast_I110_Y (.A(I110_un1_Y), .B(N428), 
        .Y(N481));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I211_un1_Y_0 (.A(N478), .B(N486)
        , .C(N493), .Y(ADD_26x26_fast_I211_un1_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I90_Y (.A(N408), .B(N412), .Y(
        N461));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I233_Y (.A(\un1_next_int[3] ), 
        .B(\integ[3]_net_1 ), .C(N491), .Y(\un1_integ[3] ));
    NOR3A inf_abs0_a_0_I_31 (.A(\DWACT_FINC_E[6] ), .B(sr_new[9]), .C(
        sr_new[10]), .Y(N_3_1));
    OA1A un1_integ_0_0_ADD_26x26_fast_I47_Y (.A(
        \un1_next_int_0_iv_0[13] ), .B(integral[14]), .C(N357), .Y(
        N415));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I119_Y (.A(N441), .B(N437), .Y(
        N490));
    MX2 \inf_abs0[7]  (.A(sr_new[7]), .B(\inf_abs0_a_0[7] ), .S(
        sr_new_1_0), .Y(\inf_abs0[7]_net_1 ));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I70_Y (.A(N320), .B(
        \integ[2]_net_1 ), .C(\un1_next_int[2] ), .Y(N438));
    DFN1E0C0 \integ[5]  (.D(\un1_integ[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(\integ[5]_net_1 ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I44_Y (.A(integral[14]), .B(
        integral[15]), .C(\un1_next_int_0_iv_0[13] ), .Y(N412));
    AX1D un1_integ_0_0_ADD_26x26_fast_I245_Y (.A(N521), .B(I188_un1_Y), 
        .C(ADD_26x26_fast_I245_Y_0), .Y(\un1_integ[15] ));
    NOR2B \state_RNICIOR2[0]  (.A(\inf_abs0[8]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[8] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I95_Y (.A(N413), .B(N417), .Y(
        N466));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y_0 (.A(\un2_next_int_m[9] )
        , .B(\un1_next_int_iv_1[9] ), .C(integral[9]), .Y(
        ADD_26x26_fast_I239_Y_0));
    DFN1E0C0 \integ[2]  (.D(\un1_integ[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(\integ[2]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I135_Y (.A(N458), .B(N466), .Y(
        N512));
    NOR3B \state_RNI3HKG3[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[11]_net_1 ), .Y(\un2_next_int_m[11] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I88_Y (.A(N410), .B(N406), .Y(
        N459));
    AX1D un1_integ_0_0_ADD_26x26_fast_I247_Y (.A(I212_un1_Y), .B(
        ADD_26x26_fast_I212_Y_0), .C(ADD_26x26_fast_I247_Y_0), .Y(
        \un1_integ[17] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I237_Y_0 (.A(\un2_next_int_m[7] )
        , .B(\un1_next_int_iv_1[7] ), .C(integral[7]), .Y(
        ADD_26x26_fast_I237_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I143_Y (.A(N466), .B(N474), .Y(
        N520));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I57_Y (.A(N345), .B(N342), .Y(
        N425));
    OA1 un1_integ_0_0_ADD_26x26_fast_I186_un1_Y (.A(N481), .B(
        I158_un1_Y), .C(N520), .Y(I186_un1_Y));
    NOR3 inf_abs0_a_0_I_29 (.A(sr_new[7]), .B(sr_new[6]), .C(sr_new[8])
        , .Y(\DWACT_FINC_E_0[5] ));
    DFN1E0C0 \integ[23]  (.D(\un1_integ[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[23]));
    OR2 un1_integ_0_0_ADD_26x26_fast_I8_P0N (.A(\un1_next_int[8] ), .B(
        integral[8]), .Y(N342));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_2 (.A(
        ADD_26x26_fast_I206_un1_Y_0), .B(N522), .C(
        ADD_26x26_fast_I206_Y_1), .Y(ADD_26x26_fast_I206_Y_2));
    AO1 un1_integ_0_0_ADD_26x26_fast_I54_Y (.A(N344), .B(N348), .C(
        N347), .Y(N422));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I131_Y (.A(N454), .B(N462), .Y(
        N508));
    XNOR2 inf_abs0_a_0_I_26 (.A(sr_new[9]), .B(N_5), .Y(
        \inf_abs0_a_0[9] ));
    NOR3B inf_abs1_a_1_I_19 (.A(\DWACT_FINC_E[2] ), .B(
        \DWACT_FINC_E_0[0] ), .C(sr_old[6]), .Y(N_7));
    NOR3B \state_RNIINCI1[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[4] ), .Y(\un2_next_int_m[4] ));
    NOR3B inf_abs1_a_1_I_16 (.A(\DWACT_FINC_E[1] ), .B(
        \DWACT_FINC_E_0[0] ), .C(sr_old[5]), .Y(N_8));
    AX1D un1_integ_0_0_ADD_26x26_fast_I254_Y (.A(I205_un1_Y), .B(
        ADD_26x26_fast_I205_Y_3), .C(ADD_26x26_fast_I254_Y_0), .Y(
        \un1_integ[24] ));
    DFN1E0C0 \integ[19]  (.D(\un1_integ[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[19]));
    NOR2 inf_abs0_a_0_I_15 (.A(sr_new[3]), .B(sr_new[4]), .Y(
        \DWACT_FINC_E_0[1] ));
    NOR2B \state_RNIR8H53[0]  (.A(\inf_abs0[10]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[10] ));
    MX2 \inf_abs1[8]  (.A(sr_old[8]), .B(\inf_abs1_a_1[8] ), .S(
        sr_old[12]), .Y(\inf_abs1[8]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I161_un1_Y (.A(N486), .B(N493), 
        .Y(I161_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I117_Y (.A(N439), .B(N435), .Y(
        N488));
    DFN1E0C0 \integ[17]  (.D(\un1_integ[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[17]));
    XOR2 inf_abs0_a_0_I_5 (.A(sr_new[0]), .B(sr_new[1]), .Y(
        \inf_abs0_a_0[1] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I33_Y (.A(integral[20]), .B(
        integral[21]), .C(\un1_next_int_0_iv[13] ), .Y(N401));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I255_Y_0 (.A(integral[25]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I255_Y_0));
    DFN1E0C0 \integ[14]  (.D(\un1_integ[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[14]));
    XNOR2 inf_abs0_a_0_I_17 (.A(sr_new[6]), .B(N_8_0), .Y(
        \inf_abs0_a_0[6] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I87_Y (.A(N409), .B(N405), .Y(
        N458));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y_0 (.A(\integ[2]_net_1 ), 
        .B(\un1_next_int[2] ), .Y(ADD_26x26_fast_I232_Y_0));
    NOR3B \state_RNIUV1L2[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[6]_net_1 ), .Y(\un2_next_int_m[6] ));
    OR3 \state_RNIT0BB1[1]  (.A(\inf_abs0_m[5] ), .B(
        \un18_next_int_m[5] ), .C(\inf_abs1_m[5] ), .Y(
        \un1_next_int_iv_1[5] ));
    MX2 \inf_abs1[0]  (.A(sr_old[0]), .B(sr_old[0]), .S(sr_old[12]), 
        .Y(\inf_abs1[0]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I84_Y (.A(N402), .B(N406), .Y(
        N455));
    MX2 \inf_abs1[11]  (.A(sr_old[11]), .B(\inf_abs1_a_1[11] ), .S(
        sr_old[12]), .Y(\inf_abs1[11]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I11_G0N (.A(\un1_next_int[11] ), 
        .B(integral[11]), .Y(N350));
    NOR2 \state_RNI5T1E[0]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 )
        , .Y(N_46_1));
    MX2 \inf_abs1[2]  (.A(sr_old[2]), .B(\inf_abs1_a_1[2] ), .S(
        sr_old[12]), .Y(\inf_abs1[2]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I140_Y (.A(N471), .B(N464), .C(
        N463), .Y(N517));
    NOR3B \state_RNIGG7R1[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[2]_net_1 ), .Y(\un2_next_int_m[2] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I149_Y (.A(N480), .B(N472), .Y(
        N526));
    OR3 \state_RNIPEN14[0]  (.A(\inf_abs0_m[2] ), .B(
        \un1_next_int_iv_0[2] ), .C(\un2_next_int_m[2] ), .Y(
        \un1_next_int[2] ));
    DFN1E0C0 \integ[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[25]));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I247_Y_0 (.A(integral[17]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I247_Y_0));
    NOR2B \state_RNIKLDA3[0]  (.A(\inf_abs0[11]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[11] ));
    MX2 \inf_abs1[6]  (.A(sr_old[6]), .B(\inf_abs1_a_1[6] ), .S(
        sr_old[12]), .Y(\inf_abs1[6]_net_1 ));
    NOR3 inf_abs0_a_0_I_33 (.A(sr_new[10]), .B(sr_new[9]), .C(
        sr_new[11]), .Y(\DWACT_FINC_E[7] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I242_Y (.A(N527), .B(I191_un1_Y), 
        .C(ADD_26x26_fast_I242_Y_0), .Y(\un1_integ[12] ));
    XNOR2 inf_abs0_a_0_I_20 (.A(sr_new[7]), .B(N_7_0), .Y(
        \inf_abs0_a_0[7] ));
    DFN1E0C0 \integ[11]  (.D(\un1_integ[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[11]));
    MX2 \inf_abs0[8]  (.A(sr_new[8]), .B(\inf_abs0_a_0[8] ), .S(
        sr_new_1_0), .Y(\inf_abs0[8]_net_1 ));
    NOR3B \state_RNIVEAE1[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[0]_net_1 ), .Y(\un2_next_int_m[0] ));
    DFN1E0C0 \integ[16]  (.D(\un1_integ[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[16]));
    XNOR2 inf_abs1_a_1_I_28 (.A(sr_old[10]), .B(N_4), .Y(
        \inf_abs1_a_1[10] ));
    NOR3 inf_abs1_a_1_I_10 (.A(sr_old[1]), .B(sr_old[0]), .C(sr_old[2])
        , .Y(\DWACT_FINC_E_0[0] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I254_Y_0 (.A(integral[24]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I254_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I163_Y (.A(I163_un1_Y), .B(N489), 
        .Y(N543));
    MX2B un1_next_int_0_sqmuxa_0__m2 (.A(sr_new_0_0), .B(sr_old[12]), 
        .S(\state[1]_net_1 ), .Y(N_3));
    AO1 un1_integ_0_0_ADD_26x26_fast_I96_Y (.A(N418), .B(N415), .C(
        N414), .Y(N467));
    MX2 \inf_abs0[10]  (.A(sr_new[10]), .B(\inf_abs0_a_0[10] ), .S(
        sr_new_1_0), .Y(\inf_abs0[10]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I114_Y (.A(I114_un1_Y), .B(N432), 
        .Y(N485));
    OA1 un1_integ_0_0_ADD_26x26_fast_I189_un1_Y (.A(N485), .B(
        I161_un1_Y), .C(N524), .Y(I189_un1_Y));
    NOR2 inf_abs0_a_0_I_21 (.A(sr_new[6]), .B(sr_new[7]), .Y(
        \DWACT_FINC_E_0[3] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I147_Y (.A(N478), .B(N470), .Y(
        N524));
    DFN1E0C0 \integ[9]  (.D(\un1_integ[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(integral[9]));
    XA1A \state_RNIQ33I[1]  (.A(sr_old[12]), .B(\inf_abs1[6]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[6] ));
    NOR2B \state_RNIONFD[1]  (.A(\inf_abs1_a_1[9] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[9] ));
    INV \integ_RNIEHQB[24]  (.A(integral[24]), .Y(integral_i[24]));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I242_Y_0 (.A(integral[12]), .B(
        \un1_next_int[12] ), .Y(ADD_26x26_fast_I242_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I235_Y (.A(N487), .B(I162_un1_Y), 
        .C(ADD_26x26_fast_I235_Y_0), .Y(\un1_integ[5] ));
    XA1A \state_RNI5I5H[1]  (.A(sr_old[12]), .B(\inf_abs1[0]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[0] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I212_Y_0 (.A(N533), .B(N518), .C(
        N517), .Y(ADD_26x26_fast_I212_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I63_Y (.A(N333), .B(N336), .Y(
        N431));
    NOR2A inf_abs1_a_1_I_11 (.A(\DWACT_FINC_E_0[0] ), .B(sr_old[3]), 
        .Y(N_10_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I118_Y (.A(I118_un1_Y), .B(N436), 
        .Y(N489));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I237_Y (.A(
        ADD_26x26_fast_I237_Y_0), .B(N537), .Y(\un1_integ[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I133_Y (.A(N464), .B(N456), .Y(
        N510));
    MX2 \inf_abs0[2]  (.A(sr_new[2]), .B(\inf_abs0_a_0[2] ), .S(
        sr_new_1_0), .Y(\inf_abs0[2]_net_1 ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I30_Y (.A(integral[21]), .B(
        integral[22]), .C(\un1_next_int_0_iv_0[13] ), .Y(N398));
    DFN1E0C0 \integ[22]  (.D(\un1_integ[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[22]));
    NOR3 inf_abs1_a_1_I_8 (.A(sr_old[1]), .B(sr_old[0]), .C(sr_old[2]), 
        .Y(N_11));
    AO1B un1_integ_0_0_ADD_26x26_fast_I43_Y (.A(integral[16]), .B(
        integral[15]), .C(\un1_next_int_0_iv_0[13] ), .Y(N411));
    DFN1E0C0 \integ_0[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral_0_0));
    OR3 un1_integ_0_0_ADD_26x26_fast_I192_Y (.A(N475), .B(I152_un1_Y), 
        .C(I192_un1_Y), .Y(N649));
    DFN1E0C0 \integ[1]  (.D(\un1_integ[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(\integ[1]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I35_Y (.A(integral[19]), .B(
        integral[20]), .C(\un1_next_int_0_iv[13] ), .Y(N403));
    NOR3B \state_RNI85UB1[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[3] ), .Y(\un2_next_int_m[3] ));
    NOR2B inf_abs0_a_0_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I53_Y (.A(N351), .B(N348), .Y(
        N421));
    AO1 un1_integ_0_0_ADD_26x26_fast_I160_Y (.A(N484), .B(N491), .C(
        N483), .Y(N537));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I91_Y (.A(N409), .B(N413), .Y(
        N462));
    AO1B un1_integ_0_0_ADD_26x26_fast_I79_Y_0 (.A(integral[23]), .B(
        integral[22]), .C(\un1_next_int_0_iv_0[13] ), .Y(
        ADD_26x26_fast_I79_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I250_Y (.A(I178_un1_Y), .B(
        ADD_26x26_fast_I209_Y_1), .C(ADD_26x26_fast_I250_Y_0), .Y(
        \un1_integ[20] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_0 (.A(N467), .B(N460), .C(
        N459), .Y(ADD_26x26_fast_I210_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I71_Y (.A(\integ[2]_net_1 ), .B(
        \un1_next_int[2] ), .C(N321), .Y(N439));
    DFN1E0C0 \integ[20]  (.D(\un1_integ[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[20]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I244_Y (.A(N523), .B(I189_un1_Y), 
        .C(ADD_26x26_fast_I244_Y_0), .Y(\un1_integ[14] ));
    NOR3 inf_abs1_a_1_I_29 (.A(sr_old[6]), .B(sr_old[8]), .C(sr_old[7])
        , .Y(\DWACT_FINC_E[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_1 (.A(N461), .B(N454), .C(
        ADD_26x26_fast_I207_Y_0), .Y(ADD_26x26_fast_I207_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I106_Y (.A(N428), .B(N425), .C(
        N424), .Y(N477));
    XNOR2 inf_abs0_a_0_I_32 (.A(sr_new[11]), .B(N_3_1), .Y(
        \inf_abs0_a_0[11] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_1 (.A(
        ADD_26x26_fast_I208_un1_Y_0), .B(N526), .C(
        ADD_26x26_fast_I208_Y_0), .Y(ADD_26x26_fast_I208_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I102_Y (.A(N424), .B(N421), .C(
        N420), .Y(N473));
    AX1D un1_integ_0_0_ADD_26x26_fast_I251_Y (.A(I176_un1_Y), .B(
        ADD_26x26_fast_I208_Y_1), .C(ADD_26x26_fast_I251_Y_0), .Y(
        \un1_integ[21] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I121_un1_Y (.A(N441), .B(
        \un1_next_int[0] ), .Y(I121_un1_Y));
    XNOR2 inf_abs1_a_1_I_26 (.A(sr_old[9]), .B(N_5_0), .Y(
        \inf_abs1_a_1[9] ));
    DFN1E0C0 \integ[18]  (.D(\un1_integ[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[18]));
    XA1A \state_RNIA58S[1]  (.A(sr_old[12]), .B(\inf_abs1[10]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[10] ));
    NOR2B \state_RNIA2CI[0]  (.A(sr_new[9]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[9] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I144_Y (.A(N475), .B(N468), .C(
        N467), .Y(N521));
    NOR3B \state_RNICMGR2[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[7]_net_1 ), .Y(\un2_next_int_m[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I83_Y (.A(N405), .B(N401), .Y(
        N454));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_0 (.A(N465), .B(N458), .C(
        N457), .Y(ADD_26x26_fast_I209_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I207_Y_0 (.A(N404), .B(N400), .Y(
        ADD_26x26_fast_I207_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I148_Y (.A(I148_un1_Y), .B(N471), 
        .Y(N525));
    NOR2B \state_RNIQMMC[1]  (.A(\inf_abs1_a_1[4] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[4] ));
    OR3 \state_RNIFIHD7[0]  (.A(\inf_abs0_m[10] ), .B(
        \un1_next_int_iv_0[10] ), .C(\un2_next_int_m[10] ), .Y(
        \un1_next_int[10] ));
    OR2 \state_RNIUVH73[1]  (.A(\un1_next_int_iv_0[7] ), .B(
        \inf_abs0_m[7] ), .Y(\un1_next_int_iv_1[7] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I60_Y (.A(N335), .B(N339), .C(
        N338), .Y(N428));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y (.A(
        ADD_26x26_fast_I232_Y_0), .B(N493), .Y(\un1_integ[2] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I204_Y_2 (.A(N398), .B(
        ADD_26x26_fast_I204_Y_0), .C(N455), .Y(ADD_26x26_fast_I204_Y_2)
        );
    NOR3B \state_RNITARO1[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[5] ), .Y(\un2_next_int_m[5] ));
    DFN1C0 \state[1]  (.D(\state_RNO_0[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[1]_net_1 ));
    XNOR2 inf_abs0_a_0_I_23 (.A(sr_new[8]), .B(N_6_0), .Y(
        \inf_abs0_a_0[8] ));
    NOR2B \state_RNIGJ381[0]  (.A(\inf_abs0[0]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[0] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I210_Y (.A(I180_un1_Y), .B(
        ADD_26x26_fast_I210_Y_0), .C(I210_un1_Y), .Y(N629));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I118_un1_Y (.A(N440), .B(N437), 
        .Y(I118_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I110_un1_Y (.A(N339), .B(N336), 
        .C(N432), .Y(I110_un1_Y));
    NOR3A inf_abs1_a_1_I_13 (.A(\DWACT_FINC_E_0[0] ), .B(sr_old[3]), 
        .C(sr_old[4]), .Y(N_9));
    MX2 \inf_abs1[7]  (.A(sr_old[7]), .B(\inf_abs1_a_1[7] ), .S(
        sr_old[12]), .Y(\inf_abs1[7]_net_1 ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I9_G0N (.A(\un2_next_int_m[9] ), 
        .B(\un1_next_int_iv_1[9] ), .C(integral[9]), .Y(N344));
    OA1B un1_integ_0_0_ADD_26x26_fast_I40_Y (.A(integral[16]), .B(
        integral[17]), .C(\un1_next_int_0_iv_0[13] ), .Y(N408));
    OA1 un1_integ_0_0_ADD_26x26_fast_I65_Y (.A(\integ[4]_net_1 ), .B(
        \un1_next_int[4] ), .C(N333), .Y(N433));
    OA1 un1_integ_0_0_ADD_26x26_fast_I207_un1_Y_0 (.A(N485), .B(
        I161_un1_Y), .C(N508), .Y(ADD_26x26_fast_I207_un1_Y_0));
    NOR2B \state_RNIF4RE2[0]  (.A(\inf_abs0[6]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[6] ));
    NOR3 inf_abs0_a_0_I_8 (.A(sr_new[1]), .B(sr_new[0]), .C(sr_new[2]), 
        .Y(N_11_0));
    AND3 inf_abs1_a_1_I_30 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E_0[6] ));
    XNOR2 inf_abs0_a_0_I_35 (.A(sr_new[12]), .B(N_2), .Y(
        \inf_abs0_a_0[12] ));
    NOR3A \state_RNIOC3C[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), .C(
        sr_old[4]), .Y(\un18_next_int_m[4] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y (.A(
        ADD_26x26_fast_I211_Y_1_0), .B(ADD_26x26_fast_I211_Y_1_tz), .C(
        ADD_26x26_fast_I211_Y_0), .Y(N631));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I178_un1_Y (.A(N512), .B(N527), 
        .Y(I178_un1_Y));
    AO1B un1_integ_0_0_ADD_26x26_fast_I45_Y (.A(integral[15]), .B(
        integral[14]), .C(\un1_next_int_0_iv_0[13] ), .Y(N413));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I137_Y (.A(N460), .B(N468), .Y(
        N514));
    XNOR2 inf_abs0_a_0_I_9 (.A(sr_new[3]), .B(N_11_0), .Y(
        \inf_abs0_a_0[3] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I3_P0N (.A(\un1_next_int[3] ), .B(
        \integ[3]_net_1 ), .Y(N327));
    NOR2B \state_RNO[0]  (.A(N_46_1), .B(calc_int), .Y(
        \state_RNO[0]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I50_Y (.A(N350), .B(N354), .C(
        N353), .Y(N418));
    AO1 un1_integ_0_0_ADD_26x26_fast_I204_Y_3 (.A(N502), .B(N517), .C(
        ADD_26x26_fast_I204_Y_2), .Y(ADD_26x26_fast_I204_Y_3));
    XNOR2 inf_abs1_a_1_I_20 (.A(sr_old[7]), .B(N_7), .Y(
        \inf_abs1_a_1[7] ));
    NOR2B \state_RNI5TBI[0]  (.A(sr_new[4]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[4] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I36_Y (.A(integral[19]), .B(
        integral[18]), .C(\un1_next_int_0_iv[13] ), .Y(N404));
    NOR2B \state_RNI6UBI[0]  (.A(sr_new[5]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[5] ));
    NOR3A inf_abs1_a_1_I_31 (.A(\DWACT_FINC_E_0[6] ), .B(sr_old[9]), 
        .C(sr_old[10]), .Y(N_3_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I0_P0N (.A(N_3), .B(
        \integ[0]_net_1 ), .Y(N318));
    NOR2 inf_abs1_a_1_I_6 (.A(sr_old[0]), .B(sr_old[1]), .Y(N_12_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I55_Y (.A(N348), .B(N345), .Y(
        N423));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I205_un1_Y (.A(N520), .B(N504), 
        .C(N658), .Y(I205_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I163_un1_Y (.A(N490), .B(
        \un1_next_int[0] ), .Y(I163_un1_Y));
    OR2 \state_RNIGQRN_0[1]  (.A(next_int_1_sqmuxa), .B(
        next_int_0_sqmuxa_1), .Y(\un1_next_int_0_iv[13] ));
    NOR2 inf_abs1_a_1_I_21 (.A(sr_old[6]), .B(sr_old[7]), .Y(
        \DWACT_FINC_E[3] ));
    OR3 \state_RNIG75G6[0]  (.A(\inf_abs0_m[8] ), .B(
        \un1_next_int_iv_0[8] ), .C(\un2_next_int_m[8] ), .Y(
        \un1_next_int[8] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I206_Y_1 (.A(N398), .B(N402), .C(
        N459), .Y(ADD_26x26_fast_I206_Y_1));
    OA1 un1_integ_0_0_ADD_26x26_fast_I5_G0N (.A(\un2_next_int_m[5] ), 
        .B(\un1_next_int_iv_1[5] ), .C(\integ[5]_net_1 ), .Y(N332));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I114_un1_Y (.A(N436), .B(N433), 
        .Y(I114_un1_Y));
    AND3 inf_abs0_a_0_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(
        \DWACT_FINC_E[4] ));
    NOR2B \state_RNI4SBI[0]  (.A(sr_new[3]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[3] ));
    DFN1E0C0 \integ[7]  (.D(\un1_integ[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(integral[7]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_2 (.A(
        ADD_26x26_fast_I207_un1_Y_0), .B(N524), .C(
        ADD_26x26_fast_I207_Y_1), .Y(ADD_26x26_fast_I207_Y_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I4_G0N (.A(\un1_next_int[4] ), 
        .B(\integ[4]_net_1 ), .Y(N329));
    NOR3A \state_RNINB3C[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), .C(
        sr_old[3]), .Y(\un18_next_int_m[3] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I195_Y (.A(N481), .B(I158_un1_Y), 
        .C(I195_un1_Y), .Y(N658));
    NOR3B \state_RNIJ2MI2[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[9] ), .Y(\un2_next_int_m[9] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I206_un1_Y_0 (.A(N506), .B(N537)
        , .Y(ADD_26x26_fast_I206_un1_Y_0));
    XNOR2 inf_abs1_a_1_I_14 (.A(sr_old[5]), .B(N_9), .Y(
        \inf_abs1_a_1[5] ));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I234_Y (.A(\un1_next_int[4] ), 
        .B(\integ[4]_net_1 ), .C(N543), .Y(\un1_integ[4] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_2 (.A(N457), .B(N450), .C(
        ADD_26x26_fast_I205_Y_1), .Y(ADD_26x26_fast_I205_Y_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I174_un1_Y (.A(N508), .B(N523), 
        .Y(I174_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I162_un1_Y (.A(N488), .B(N442), 
        .Y(I162_un1_Y));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I240_Y (.A(\un1_next_int[10] ), 
        .B(integral[10]), .C(N652), .Y(\un1_integ[10] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I156_Y (.A(N487), .B(N480), .C(
        N479), .Y(N533));
    DFN1E0C0 \integ[8]  (.D(\un1_integ[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1), .Q(integral[8]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I85_Y (.A(N407), .B(N403), .Y(
        N456));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I251_Y_0 (.A(integral[21]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I251_Y_0));
    AND3 inf_abs0_a_0_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(N_6_0));
    OR3 un1_integ_0_0_ADD_26x26_fast_I9_P0N (.A(\un2_next_int_m[9] ), 
        .B(\un1_next_int_iv_1[9] ), .C(integral[9]), .Y(N345));
    OA1 un1_integ_0_0_ADD_26x26_fast_I208_un1_Y_0 (.A(N487), .B(
        I162_un1_Y), .C(N510), .Y(ADD_26x26_fast_I208_un1_Y_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I31_Y (.A(integral[22]), .B(
        integral[21]), .C(\un1_next_int_0_iv_0[13] ), .Y(N399));
    XNOR2 inf_abs1_a_1_I_12 (.A(sr_old[4]), .B(N_10_0), .Y(
        \inf_abs1_a_1[4] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I235_Y_0 (.A(\un2_next_int_m[5] )
        , .B(\un1_next_int_iv_1[5] ), .C(\integ[5]_net_1 ), .Y(
        ADD_26x26_fast_I235_Y_0));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I241_Y (.A(\un1_next_int[11] ), 
        .B(integral[11]), .C(N649), .Y(\un1_integ[11] ));
    NOR3 inf_abs0_a_0_I_18 (.A(sr_new[4]), .B(sr_new[3]), .C(sr_new[5])
        , .Y(\DWACT_FINC_E_0[2] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I11_P0N (.A(\un1_next_int[11] ), 
        .B(integral[11]), .Y(N351));
    NOR2B \state_RNI1L0L1[0]  (.A(\inf_abs0[2]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[2] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I243_Y_0 (.A(integral[13]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I243_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I105_Y (.A(N339), .B(N342), .C(
        N423), .Y(N476));
    MX2 \inf_abs0[11]  (.A(sr_new[11]), .B(\inf_abs0_a_0[11] ), .S(
        sr_new_1_0), .Y(\inf_abs0[11]_net_1 ));
    XOR2 inf_abs1_a_1_I_5 (.A(sr_old[0]), .B(sr_old[1]), .Y(
        \inf_abs1_a_1[1] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I101_Y (.A(N419), .B(N423), .Y(
        N472));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I66_Y (.A(N326), .B(
        \integ[4]_net_1 ), .C(\un1_next_int[4] ), .Y(N434));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I248_Y (.A(
        \un1_next_int_0_iv_0[13] ), .B(integral[18]), .C(N631), .Y(
        \un1_integ[18] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I99_Y (.A(N417), .B(N421), .Y(
        N470));
    OR2 un1_integ_0_0_ADD_26x26_fast_I92_Y (.A(N410), .B(N414), .Y(
        N463));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I191_un1_Y (.A(N528), .B(N543), 
        .Y(I191_un1_Y));
    NOR3A \state_RNIL93C[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), .C(
        sr_old[1]), .Y(\un18_next_int_m[1] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I79_Y (.A(
        ADD_26x26_fast_I79_Y_0), .B(N401), .Y(N450));
    AO1 un1_integ_0_0_ADD_26x26_fast_I72_Y (.A(N317), .B(N321), .C(
        N320), .Y(N440));
    OR2A un1_integ_0_0_ADD_26x26_fast_I13_P0N (.A(
        \un1_next_int_0_iv[13] ), .B(integral[13]), .Y(N357));
    OA1B un1_integ_0_0_ADD_26x26_fast_I46_Y (.A(integral[13]), .B(
        integral[14]), .C(\un1_next_int_0_iv_0[13] ), .Y(N414));
    NOR2B \state_RNITQ9L2[0]  (.A(\inf_abs0[7]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[7] ));
    OR2 \state_RNI98U03[1]  (.A(\un1_next_int_iv_0[6] ), .B(
        \inf_abs0_m[6] ), .Y(\un1_next_int_iv_1[6] ));
    OR3 \state_RNIVBVB1[1]  (.A(\inf_abs0_m[9] ), .B(
        \un18_next_int_m[9] ), .C(\inf_abs1_m[9] ), .Y(
        \un1_next_int_iv_1[9] ));
    NOR3 inf_abs1_a_1_I_33 (.A(sr_old[10]), .B(sr_old[9]), .C(
        sr_old[11]), .Y(\DWACT_FINC_E_0[7] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I116_Y (.A(N438), .B(N435), .C(
        N434), .Y(N487));
    AO1 un1_integ_0_0_ADD_26x26_fast_I112_Y (.A(N434), .B(N431), .C(
        N430), .Y(N483));
    NOR2A inf_abs0_a_0_I_25 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .Y(
        N_5));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I8_G0N (.A(\un1_next_int[8] ), 
        .B(integral[8]), .Y(N341));
    OR3 un1_integ_0_0_ADD_26x26_fast_I211_Y_1_tz (.A(N477), .B(
        I154_un1_Y), .C(ADD_26x26_fast_I211_un1_Y_0), .Y(
        ADD_26x26_fast_I211_Y_1_tz));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I213_un1_Y_0 (.A(N482), .B(N490)
        , .C(\un1_next_int[0] ), .Y(ADD_26x26_fast_I213_un1_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I210_un1_Y (.A(N514), .B(N491), 
        .C(N530), .Y(I210_un1_Y));
    OR2 \state_RNI780M5[0]  (.A(\un1_next_int_iv_1[6] ), .B(
        \un2_next_int_m[6] ), .Y(\un1_next_int[6] ));
    NOR3A inf_abs0_a_0_I_27 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .C(
        sr_new[9]), .Y(N_4_0));
    
endmodule


module error_calc_13s_12s_4(
       cur_error,
       LED_12_i_0,
       LED_12,
       average,
       calc_error,
       n_rst_c,
       clk_c
    );
output [12:0] cur_error;
input  LED_12_i_0;
input  [7:0] LED_12;
input  [6:2] average;
input  calc_error;
input  n_rst_c;
input  clk_c;

    wire N_38, N_40, GND, VCC;
    
    AX1B un2_diffreg_1_m37 (.A(LED_12[5]), .B(LED_12[6]), .C(LED_12[7])
        , .Y(N_38));
    DFN1E1C0 \diffreg[3]  (.D(average[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[3]));
    XNOR2 un2_diffreg_1_m39 (.A(LED_12[6]), .B(LED_12[5]), .Y(N_40));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \diffreg[7]  (.D(LED_12[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[7]));
    DFN1E1C0 \diffreg[1]  (.D(average[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[1]));
    DFN1E1C0 \diffreg[12]  (.D(N_38), .CLK(clk_c), .CLR(n_rst_c), .E(
        calc_error), .Q(cur_error[12]));
    DFN1E1C0 \diffreg[11]  (.D(N_40), .CLK(clk_c), .CLR(n_rst_c), .E(
        calc_error), .Q(cur_error[11]));
    GND GND_i (.Y(GND));
    DFN1E1C0 \diffreg[9]  (.D(LED_12[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[9]));
    DFN1E1C0 \diffreg[8]  (.D(LED_12[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[8]));
    DFN1E1C0 \diffreg[6]  (.D(LED_12[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[6]));
    DFN1E1C0 \diffreg[10]  (.D(LED_12_i_0), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[10]));
    DFN1E1C0 \diffreg[5]  (.D(LED_12[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[5]));
    DFN1E1C0 \diffreg[4]  (.D(average[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[4]));
    DFN1E1C0 \diffreg[2]  (.D(average[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[2]));
    DFN1E1C0 \diffreg[0]  (.D(average[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[0]));
    
endmodule


module derivative_calc_13s_4(
       derivative_0,
       sr_prev,
       sr_new,
       sr_new_0_0,
       deriv_enable,
       n_rst_c,
       clk_c
    );
output derivative_0;
input  [12:0] sr_prev;
input  [11:0] sr_new;
input  sr_new_0_0;
input  deriv_enable;
input  n_rst_c;
input  clk_c;

    wire SUB_13x13_medium_area_I49_Y_1, N208, N176, 
        SUB_13x13_medium_area_I49_Y_0, 
        SUB_13x13_medium_area_I26_un1_Y_0, 
        SUB_13x13_medium_area_I49_un1_Y_1, 
        SUB_13x13_medium_area_I49_un1_Y_0, N_15, 
        SUB_13x13_medium_area_I42_Y_1, N218, N180, 
        SUB_13x13_medium_area_I42_Y_0, 
        SUB_13x13_medium_area_I30_un1_Y_0, 
        SUB_13x13_medium_area_I42_un1_Y_1, N_9, N_7, 
        SUB_13x13_medium_area_I41_Y_0, 
        SUB_13x13_medium_area_I34_un1_Y_0, 
        SUB_13x13_medium_area_I41_un1_Y_0, N_5, 
        SUB_13x13_medium_area_I28_un1_Y_0, 
        SUB_13x13_medium_area_I32_un1_Y_0, N_24, N226, N204, N212, 
        N222, N185, N_21, N_13, GND, VCC;
    
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I34_un1_Y_0 (.A(
        sr_new[1]), .B(sr_prev[1]), .Y(
        SUB_13x13_medium_area_I34_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y_0 (.A(
        SUB_13x13_medium_area_I30_un1_Y_0), .B(sr_new[6]), .C(
        sr_prev[6]), .Y(SUB_13x13_medium_area_I42_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I15_S (.A(sr_prev[2]), 
        .B(sr_new[2]), .Y(N_5));
    OR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I36_Y (.A(sr_prev[0]), 
        .B(sr_new[0]), .Y(N185));
    XNOR3 un2_deriv_out_0_0_SUB_13x13_medium_area_I82_Y (.A(sr_new_0_0)
        , .B(sr_prev[12]), .C(N226), .Y(N_24));
    VCC VCC_i (.Y(VCC));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I64_Y (.A(N204), .B(
        sr_new[11]), .C(sr_prev[11]), .Y(N226));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I41_Y_0 (.A(
        SUB_13x13_medium_area_I34_un1_Y_0), .B(sr_new[2]), .C(
        sr_prev[2]), .Y(SUB_13x13_medium_area_I41_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I19_S (.A(sr_prev[6]), 
        .B(sr_new[6]), .Y(N_13));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I28_Y (.A(
        SUB_13x13_medium_area_I28_un1_Y_0), .B(sr_new[8]), .C(
        sr_prev[8]), .Y(N208));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y_1 (.A(N218), .B(
        N180), .C(SUB_13x13_medium_area_I42_Y_0), .Y(
        SUB_13x13_medium_area_I42_Y_1));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I28_un1_Y_0 (.A(
        sr_new[7]), .B(sr_prev[7]), .Y(
        SUB_13x13_medium_area_I28_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y_0 (.A(
        SUB_13x13_medium_area_I26_un1_Y_0), .B(sr_new[10]), .C(
        sr_prev[10]), .Y(SUB_13x13_medium_area_I49_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I20_S (.A(sr_prev[7]), 
        .B(sr_new[7]), .Y(N_15));
    DFN1E1C0 \deriv_out[12]  (.D(N_24), .CLK(clk_c), .CLR(n_rst_c), .E(
        deriv_enable), .Q(derivative_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I17_S (.A(sr_prev[4]), 
        .B(sr_new[4]), .Y(N_9));
    GND GND_i (.Y(GND));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I23_S (.A(sr_prev[10])
        , .B(sr_new[10]), .Y(N_21));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I26_un1_Y_0 (.A(
        sr_new[9]), .B(sr_prev[9]), .Y(
        SUB_13x13_medium_area_I26_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I32_Y (.A(
        SUB_13x13_medium_area_I32_un1_Y_0), .B(sr_new[4]), .C(
        sr_prev[4]), .Y(N218));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I30_un1_Y_0 (.A(
        sr_new[5]), .B(sr_prev[5]), .Y(
        SUB_13x13_medium_area_I30_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y (.A(
        SUB_13x13_medium_area_I49_un1_Y_1), .B(N212), .C(
        SUB_13x13_medium_area_I49_Y_1), .Y(N204));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I32_un1_Y_0 (.A(
        sr_new[3]), .B(sr_prev[3]), .Y(
        SUB_13x13_medium_area_I32_un1_Y_0));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I31_Y (.A(sr_new[5]), 
        .B(sr_prev[5]), .C(N_13), .Y(N180));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I41_un1_Y_0 (.A(
        sr_new[1]), .B(sr_prev[1]), .C(N_5), .Y(
        SUB_13x13_medium_area_I41_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y_1 (.A(N208), .B(
        N176), .C(SUB_13x13_medium_area_I49_Y_0), .Y(
        SUB_13x13_medium_area_I49_Y_1));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I16_S (.A(sr_prev[3]), 
        .B(sr_new[3]), .Y(N_7));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y (.A(
        SUB_13x13_medium_area_I42_un1_Y_1), .B(N222), .C(
        SUB_13x13_medium_area_I42_Y_1), .Y(N212));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I27_Y (.A(sr_new[9]), 
        .B(sr_prev[9]), .C(N_21), .Y(N176));
    NOR2B un2_deriv_out_0_0_SUB_13x13_medium_area_I49_un1_Y_1 (.A(
        SUB_13x13_medium_area_I49_un1_Y_0), .B(N176), .Y(
        SUB_13x13_medium_area_I49_un1_Y_1));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I49_un1_Y_0 (.A(
        sr_new[8]), .B(sr_prev[8]), .C(N_15), .Y(
        SUB_13x13_medium_area_I49_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I41_Y (.A(
        SUB_13x13_medium_area_I41_un1_Y_0), .B(N185), .C(
        SUB_13x13_medium_area_I41_Y_0), .Y(N222));
    NOR3A un2_deriv_out_0_0_SUB_13x13_medium_area_I42_un1_Y_1 (.A(N180)
        , .B(N_9), .C(N_7), .Y(SUB_13x13_medium_area_I42_un1_Y_1));
    
endmodule


module pwm_tx_200s_32s_13s_10_216s_51s(
       off_div,
       act_ctl_5_i,
       act_ctl_5_0,
       act_ctl_5_8,
       pwm_chg,
       pwm_chg_0,
       n_rst_c,
       clk_c,
       act_ctl_5,
       act_ctl_5_9,
       act_ctl_5_4,
       act_ctl_5_3,
       act_ctl_5_7,
       primary_12_c
    );
input  [31:0] off_div;
input  act_ctl_5_i;
input  act_ctl_5_0;
input  act_ctl_5_8;
input  pwm_chg;
input  pwm_chg_0;
input  n_rst_c;
input  clk_c;
input  act_ctl_5;
input  act_ctl_5_9;
input  act_ctl_5_4;
input  act_ctl_5_3;
input  act_ctl_5_7;
output primary_12_c;

    wire counter_N_3_0, I_140_0, I_140, \DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] , \DWACT_COMP0_E[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] , N_21, \counter[9]_net_1 , 
        I_6, \DWACT_FDEC_E[0] , N_5, N_17, N_13, \counter[8]_net_1 , 
        N_7, N_3, \counter[3]_net_1 , counter_m6_0_a2_7, 
        counter_m6_0_a2_2, counter_m6_0_a2_1, counter_m6_0_a2_6, 
        \counter[16]_net_1 , \counter[18]_net_1 , counter_m6_0_a2_4, 
        \counter[15]_net_1 , \counter[10]_net_1 , \counter[17]_net_1 , 
        \counter[13]_net_1 , \counter[14]_net_1 , \counter[11]_net_1 , 
        \counter[12]_net_1 , \counter_RNO[1]_net_1 , counter_N_8_0, 
        \counter_RNO_1[1]_net_1 , counter_N_7_0, counter_c18, 
        counter_c8, cur_pwm_RNO_net_1, \counter[1]_net_1 , 
        \counter[0]_net_1 , \counter_RNO[0]_net_1 , d_N_3_mux_4, 
        counter_N_3_mux, counter_N_7, \counter_RNO_0[31]_net_1 , 
        \counter[31]_net_1 , \counter[30]_net_1 , counter_c29, 
        cur_pwm_RNIA74H44_0_net_1, counter_n30, counter_n29, 
        \counter[29]_net_1 , counter_c28, counter_n28, counter_n28_tz, 
        \counter[27]_net_1 , counter_c26, \counter[28]_net_1 , 
        counter_n27, counter_n26, counter_n26_tz, \counter[25]_net_1 , 
        counter_c24, \counter[26]_net_1 , counter_n25, counter_n24, 
        counter_n24_tz, \counter[23]_net_1 , counter_c22, 
        \counter[24]_net_1 , counter_n23, counter_n22, counter_n22_tz, 
        \counter[21]_net_1 , counter_c20, \counter[22]_net_1 , 
        counter_n21, counter_n20, counter_n20_tz, \counter[19]_net_1 , 
        \counter[20]_net_1 , counter_n19, counter_n18, counter_c17, 
        counter_n17, counter_c16, counter_n16, counter_c15, 
        counter_n15, counter_c14, counter_n14, counter_c13, 
        counter_n13, counter_c12, counter_n12, counter_c11, 
        counter_n11, counter_c10, counter_n10, counter_n10_tz, 
        counter_n9, counter_n8, counter_n8_tz, \counter[7]_net_1 , 
        counter_c6, counter_n7, counter_n6, counter_n6_tz, 
        \counter[5]_net_1 , counter_c4, \counter[6]_net_1 , counter_n5, 
        counter_n4, counter_n4_tz, counter_c2, \counter[4]_net_1 , 
        counter_n3, counter_n2, counter_n2_tz, \counter[2]_net_1 , 
        \off_time[2] , \off_reg[2]_net_1 , \off_time[8] , 
        \off_reg[8]_net_1 , \off_time[9] , \off_reg[9]_net_1 , 
        \off_time[10] , \off_reg[10]_net_1 , \off_time[11] , 
        \off_reg[11]_net_1 , \off_time[12] , \off_reg[12]_net_1 , 
        \off_time[13] , \off_reg[13]_net_1 , \off_time[20] , 
        \off_reg[20]_net_1 , \off_time[6] , \off_reg[6]_net_1 , 
        \off_time[1] , \off_reg[1]_net_1 , \off_time[0] , 
        \off_reg[0]_net_1 , \off_time[4] , \off_reg[4]_net_1 , 
        \off_time[7] , \off_reg[7]_net_1 , \off_time[18] , 
        \off_reg[18]_net_1 , \off_time[22] , \off_reg[22]_net_1 , 
        \off_time[24] , \off_reg[24]_net_1 , \off_time[25] , 
        \off_reg[25]_net_1 , \off_time[26] , \off_reg[26]_net_1 , 
        \off_time[23] , \off_reg[23]_net_1 , \off_time[28] , 
        \off_reg[28]_net_1 , \off_time[21] , \off_reg[21]_net_1 , 
        \off_time[29] , \off_reg[29]_net_1 , \off_time[27] , 
        \off_reg[27]_net_1 , \off_time[14] , \off_reg[14]_net_1 , 
        \off_time[15] , \off_reg[15]_net_1 , \off_time[3] , 
        \off_reg[3]_net_1 , \off_time[31] , \off_reg[31]_net_1 , 
        \off_time[5] , \off_reg[5]_net_1 , \off_time[30] , 
        \off_reg[30]_net_1 , \off_time[19] , \off_reg[19]_net_1 , 
        \off_time[17] , \off_reg[17]_net_1 , \off_time[16] , 
        \off_reg[16]_net_1 , \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] , N_11, N_10, N_9, N_6, 
        N_8, I_12_0, N_16, N_18, I_20_0, N_12, I_17_0, N_14, I_14_0, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] , \DWACT_BL_EQUAL_0_E[0] , 
        \DWACT_BL_EQUAL_0_E[1] , \DWACT_BL_EQUAL_0_E[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] , \DWACT_COMP0_E_0[1] , 
        \DWACT_COMP0_E_0[2] , \DWACT_COMP0_E[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] , N_11_0, N_10_0, N_9_0, 
        N_6_0, N_8_0, N_7_0, N_5_0, N_2, N_3_0, N_4, N_21_0, N_20, 
        N_19, N_16_0, N_18_0, N_17_0, N_15, N_12_0, N_13_0, N_14_0, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] , 
        \DWACT_BL_EQUAL_0_E[4] , \DWACT_BL_EQUAL_0_E[3] , 
        \DWACT_BL_EQUAL_0_E_0[0] , \DWACT_BL_EQUAL_0_E_0[1] , 
        \DWACT_BL_EQUAL_0_E_0[2] , \DWACT_CMPLE_PO0_DWACT_COMP0_E[1] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[0] , N_31, N_30, N_29, N_26, 
        N_28, N_27, N_25, N_22, N_23, N_24, \ACT_LT4_E[3] , 
        \ACT_LT4_E[6] , \ACT_LT4_E[10] , \ACT_LT4_E[7] , 
        \ACT_LT4_E[8] , \ACT_LT4_E[5] , \ACT_LT4_E[4] , \ACT_LT4_E[0] , 
        \ACT_LT4_E[1] , \ACT_LT4_E[2] , \DWACT_BL_EQUAL_0_E_0[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] , 
        \DWACT_BL_EQUAL_0_E_1[0] , \DWACT_BL_EQUAL_0_E_1[1] , 
        \DWACT_BL_EQUAL_0_E_1[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] , 
        \DWACT_BL_EQUAL_0_E_2[0] , \DWACT_BL_EQUAL_0_E_2[1] , 
        \DWACT_BL_EQUAL_0_E_2[2] , \DWACT_BL_EQUAL_0_E_1[3] , 
        \DWACT_BL_EQUAL_0_E_0[4] , \DWACT_BL_EQUAL_0_E[5] , 
        \DWACT_BL_EQUAL_0_E[6] , \DWACT_BL_EQUAL_0_E[7] , 
        \DWACT_BL_EQUAL_0_E[8] , \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] , N_41, N_40, N_39, N_36, 
        N_38, N_37, N_35, N_32, N_33, N_34, \ACT_LT3_E[3] , 
        \ACT_LT3_E[4] , \ACT_LT3_E[5] , \ACT_LT3_E[0] , \ACT_LT3_E[1] , 
        \ACT_LT3_E[2] , \DWACT_BL_EQUAL_0_E_3[2] , 
        \DWACT_BL_EQUAL_0_E_3[1] , \DWACT_BL_EQUAL_0_E_3[0] , N_51, 
        N_50, N_49, N_46, N_48, N_47, N_45, N_42, N_43, N_44, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] , 
        \DWACT_BL_EQUAL_0_E_1[4] , \DWACT_BL_EQUAL_0_E_2[3] , 
        \DWACT_BL_EQUAL_0_E_4[0] , \DWACT_BL_EQUAL_0_E_4[1] , 
        \DWACT_BL_EQUAL_0_E_4[2] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] , 
        \DWACT_BL_EQUAL_0_E[12] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] , 
        \DWACT_BL_EQUAL_0_E_5[0] , \DWACT_BL_EQUAL_0_E_5[1] , 
        \DWACT_BL_EQUAL_0_E_5[2] , \DWACT_BL_EQUAL_0_E_3[3] , 
        \DWACT_BL_EQUAL_0_E_2[4] , \DWACT_BL_EQUAL_0_E_0[5] , 
        \DWACT_BL_EQUAL_0_E_0[6] , \DWACT_BL_EQUAL_0_E_0[7] , 
        \DWACT_BL_EQUAL_0_E_0[8] , \DWACT_BL_EQUAL_0_E[9] , 
        \DWACT_BL_EQUAL_0_E[10] , \DWACT_BL_EQUAL_0_E[11] , N_2_0, 
        \DWACT_FDEC_E[2] , N_3_1, \DWACT_FDEC_E[1] , N_4_0, GND, VCC;
    
    DFN1C0 \counter[19]  (.D(counter_n19), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[19]_net_1 ));
    AND3 un1_counter_0_I_78 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] ));
    NOR2A \off_reg_RNILOVP[11]  (.A(\off_reg[11]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[11] ));
    NOR3 un1_counter_2_0_I_17 (.A(\counter[20]_net_1 ), .B(
        \counter[19]_net_1 ), .C(\counter[21]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] ));
    NOR2A \off_reg_RNIMPVP[12]  (.A(\off_reg[12]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[12] ));
    AND2A un1_counter_0_I_51 (.A(\off_time[26] ), .B(
        \counter[26]_net_1 ), .Y(\ACT_LT3_E[5] ));
    NOR2A \off_reg_RNI54FT[28]  (.A(\off_reg[28]_net_1 ), .B(act_ctl_5)
        , .Y(\off_time[28] ));
    DFN1E1C0 \off_reg[28]  (.D(off_div[28]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[28]_net_1 ));
    AX1C \counter_RNO_0[2]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .C(\counter[2]_net_1 ), .Y(counter_n2_tz));
    DFN1C0 \counter[28]  (.D(counter_n28), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[28]_net_1 ));
    XNOR2 un1_counter_0_I_73 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .Y(\DWACT_BL_EQUAL_0_E_2[2] ));
    OA1A un1_counter_0_I_136 (.A(N_6_0), .B(N_8_0), .C(N_7_0), .Y(
        N_11_0));
    OR2A un1_counter_2_0_I_116 (.A(I_17_0), .B(\counter[6]_net_1 ), .Y(
        N_12));
    OA1A un1_counter_0_I_132 (.A(\counter[3]_net_1 ), .B(\off_time[3] )
        , .C(N_3_0), .Y(N_7_0));
    DFN1E1C0 \off_reg[15]  (.D(off_div[15]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[15]_net_1 ));
    DFN1E1C0 \off_reg[26]  (.D(off_div[26]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[26]_net_1 ));
    AND3 un1_counter_0_I_14 (.A(\DWACT_BL_EQUAL_0_E[9] ), .B(
        \DWACT_BL_EQUAL_0_E[10] ), .C(\DWACT_BL_EQUAL_0_E[11] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] ));
    XA1B \counter_RNO[11]  (.A(\counter[11]_net_1 ), .B(counter_c10), 
        .C(counter_N_3_0), .Y(counter_n11));
    DFN1C0 \counter[29]  (.D(counter_n29), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[29]_net_1 ));
    DFN1E1C0 \off_reg[5]  (.D(off_div[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[5]_net_1 ));
    NOR3 un1_counter_2_0_I_77 (.A(\counter[12]_net_1 ), .B(
        \counter[10]_net_1 ), .C(\counter[11]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] ));
    XNOR2 un1_counter_0_I_82 (.A(\counter[15]_net_1 ), .B(
        \off_time[15] ), .Y(\DWACT_BL_EQUAL_0_E_1[0] ));
    DFN1C0 \counter[11]  (.D(counter_n11), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[11]_net_1 ));
    XNOR2 un1_counter_0_I_109 (.A(\counter[6]_net_1 ), .B(
        \off_time[6] ), .Y(\DWACT_BL_EQUAL_0_E_0[1] ));
    NOR2A un1_counter_2_0_I_118 (.A(I_14_0), .B(\counter[5]_net_1 ), 
        .Y(N_14));
    OR2A un1_counter_0_I_103 (.A(\counter[14]_net_1 ), .B(
        \off_time[14] ), .Y(N_29));
    NOR2A \counter_RNO[28]  (.A(counter_n28_tz), .B(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n28));
    XA1B \counter_RNO[15]  (.A(\counter[15]_net_1 ), .B(counter_c14), 
        .C(counter_N_3_0), .Y(counter_n15));
    XNOR2 un1_counter_0_I_25 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .Y(\DWACT_BL_EQUAL_0_E_2[3] ));
    AND2 un1_counter_0_I_114 (.A(\DWACT_BL_EQUAL_0_E[4] ), .B(
        \DWACT_BL_EQUAL_0_E[3] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] ));
    NOR2B \counter_RNIJR5M6[13]  (.A(counter_c12), .B(
        \counter[13]_net_1 ), .Y(counter_c13));
    XNOR2 un1_counter_0_I_11 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .Y(\DWACT_BL_EQUAL_0_E_3[3] ));
    NOR3C \counter_RNIMJ974[8]  (.A(\counter[7]_net_1 ), .B(counter_c6)
        , .C(\counter[8]_net_1 ), .Y(counter_c8));
    AX1C \counter_RNO_0[22]  (.A(\counter[21]_net_1 ), .B(counter_c20), 
        .C(\counter[22]_net_1 ), .Y(counter_n22_tz));
    NOR2A \off_reg_RNIUTFT[30]  (.A(\off_reg[30]_net_1 ), .B(act_ctl_5)
        , .Y(\off_time[30] ));
    XA1B \counter_RNO[7]  (.A(\counter[7]_net_1 ), .B(counter_c6), .C(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n7));
    OA1A un1_counter_2_0_I_125 (.A(N_16), .B(N_18), .C(N_17), .Y(N_21));
    DFN1E1C0 \off_reg[2]  (.D(off_div[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[2]_net_1 ));
    XNOR2 un1_counter_0_I_72 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .Y(\DWACT_BL_EQUAL_0_E_1[3] ));
    OA1 un1_counter_0_I_126 (.A(N_21_0), .B(N_20), .C(N_19), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] ));
    NOR2A \off_reg_RNI43FT[27]  (.A(\off_reg[27]_net_1 ), .B(act_ctl_5)
        , .Y(\off_time[27] ));
    NOR2A \off_reg_RNINQVP[13]  (.A(\off_reg[13]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[13] ));
    DFN1C0 \counter[6]  (.D(counter_n6), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[6]_net_1 ));
    AO1C un1_counter_0_I_122 (.A(\counter[7]_net_1 ), .B(\off_time[7] )
        , .C(N_12_0), .Y(N_18_0));
    NOR3C \counter_RNIDDU5D[26]  (.A(\counter[25]_net_1 ), .B(
        counter_c24), .C(\counter[26]_net_1 ), .Y(counter_c26));
    XA1B \counter_RNO[31]  (.A(\counter_RNO_0[31]_net_1 ), .B(
        \counter[31]_net_1 ), .C(counter_N_3_0), .Y(counter_N_7));
    NOR3C \counter_RNIPBQF2[18]  (.A(\counter[16]_net_1 ), .B(
        \counter[18]_net_1 ), .C(counter_m6_0_a2_4), .Y(
        counter_m6_0_a2_6));
    NOR2 un1_act_ctl_I_6 (.A(act_ctl_5_7), .B(act_ctl_5_7), .Y(I_6));
    DFN1C0 \counter[21]  (.D(counter_n21), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[21]_net_1 ));
    AND2 un1_counter_0_I_20 (.A(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] ), .B(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] ), .Y(
        \DWACT_COMP0_E_0[1] ));
    OR2 un1_act_ctl_I_10 (.A(act_ctl_5_3), .B(act_ctl_5_3), .Y(
        \DWACT_FDEC_E[0] ));
    XNOR2 un1_counter_2_0_I_109 (.A(\counter[6]_net_1 ), .B(I_17_0), 
        .Y(\DWACT_BL_EQUAL_0_E[1] ));
    XNOR2 \counter_RNO_1[1]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(\counter_RNO_1[1]_net_1 ));
    DFN1C0 \counter[3]  (.D(counter_n3), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[3]_net_1 ));
    DFN1C0 \counter[2]  (.D(counter_n2), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[2]_net_1 ));
    AND3 un1_counter_0_I_45 (.A(\DWACT_BL_EQUAL_0_E_3[2] ), .B(
        \DWACT_BL_EQUAL_0_E_3[1] ), .C(\DWACT_BL_EQUAL_0_E_3[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] ));
    DFN1E1C0 \off_reg[23]  (.D(off_div[23]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[23]_net_1 ));
    NOR2A \counter_RNO[8]  (.A(counter_n8_tz), .B(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n8));
    NOR2A un1_counter_2_0_I_121 (.A(N_13), .B(\counter[8]_net_1 ), .Y(
        N_17));
    XA1B \counter_RNO[13]  (.A(\counter[13]_net_1 ), .B(counter_c12), 
        .C(counter_N_3_0), .Y(counter_n13));
    AO1C un1_counter_0_I_57 (.A(\off_time[20] ), .B(
        \counter[20]_net_1 ), .C(N_34), .Y(N_36));
    NOR3C \counter_RNIFGLF4[11]  (.A(counter_m6_0_a2_2), .B(
        counter_m6_0_a2_1), .C(counter_m6_0_a2_6), .Y(
        counter_m6_0_a2_7));
    NOR2A \off_reg_RNI65FT[29]  (.A(\off_reg[29]_net_1 ), .B(act_ctl_5)
        , .Y(\off_time[29] ));
    DFN1E1C0 \off_reg[9]  (.D(off_div[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[9]_net_1 ));
    XNOR2 un1_counter_0_I_26 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(\DWACT_BL_EQUAL_0_E_4[2] ));
    AX1C \counter_RNO_0[4]  (.A(\counter[3]_net_1 ), .B(counter_c2), 
        .C(\counter[4]_net_1 ), .Y(counter_n4_tz));
    AO1C un1_counter_0_I_35 (.A(\off_time[28] ), .B(
        \counter[28]_net_1 ), .C(N_44), .Y(N_46));
    AO1 un1_counter_0_I_65 (.A(\DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] ), 
        .B(\DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] ), .C(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] ), .Y(\DWACT_COMP0_E[0] ));
    OR2A un1_act_ctl_I_11 (.A(act_ctl_5_3), .B(\DWACT_FDEC_E[0] ), .Y(
        N_5));
    NOR2A \off_reg_RNIPT0Q[24]  (.A(\off_reg[24]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[24] ));
    NOR2A \off_reg_RNIKNVP[10]  (.A(\off_reg[10]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[10] ));
    AND2 un1_counter_0_I_84 (.A(\DWACT_BL_EQUAL_0_E_0[3] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[1] ));
    NOR2A \off_reg_RNIVOT6[1]  (.A(\off_reg[1]_net_1 ), .B(act_ctl_5_4)
        , .Y(\off_time[1] ));
    NOR2A \off_reg_RNI0QT6[2]  (.A(\off_reg[2]_net_1 ), .B(act_ctl_5_4)
        , .Y(\off_time[2] ));
    DFN1C0 cur_pwm (.D(cur_pwm_RNO_net_1), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(primary_12_c));
    XA1B \counter_RNO[12]  (.A(\counter[12]_net_1 ), .B(counter_c11), 
        .C(counter_N_3_0), .Y(counter_n12));
    AOI1A un1_counter_0_I_95 (.A(\ACT_LT4_E[3] ), .B(\ACT_LT4_E[6] ), 
        .C(\ACT_LT4_E[10] ), .Y(\DWACT_CMPLE_PO0_DWACT_COMP0_E[0] ));
    OA1A un1_counter_0_I_40 (.A(N_46), .B(N_48), .C(N_47), .Y(N_51));
    NOR3 \counter_RNO[1]  (.A(counter_N_8_0), .B(
        \counter_RNO_1[1]_net_1 ), .C(counter_N_7_0), .Y(
        \counter_RNO[1]_net_1 ));
    DFN1C0 \counter[17]  (.D(counter_n17), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[17]_net_1 ));
    NOR2 \counter_RNO_0[1]  (.A(primary_12_c), .B(I_140_0), .Y(
        counter_N_8_0));
    OR2 un1_counter_2_0_I_129 (.A(\counter[0]_net_1 ), .B(act_ctl_5_8), 
        .Y(N_6));
    DFN1C0 \counter[4]  (.D(counter_n4), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[4]_net_1 ));
    NOR2B \counter_RNI2I3M7[15]  (.A(counter_c14), .B(
        \counter[15]_net_1 ), .Y(counter_c15));
    AND2 un1_counter_0_I_30 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] ));
    OR2A un1_counter_0_I_60 (.A(\counter[23]_net_1 ), .B(
        \off_time[23] ), .Y(N_39));
    DFN1E1C0 \off_reg[11]  (.D(off_div[11]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[11]_net_1 ));
    AND2 un1_counter_0_I_29 (.A(\DWACT_BL_EQUAL_0_E_1[4] ), .B(
        \DWACT_BL_EQUAL_0_E_2[3] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] ));
    NOR2A \off_reg_RNIT00Q[19]  (.A(\off_reg[19]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[19] ));
    DFN1E1C0 \off_reg[22]  (.D(off_div[22]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[22]_net_1 ));
    DFN1C0 \counter[10]  (.D(counter_n10), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[10]_net_1 ));
    NOR3C \counter_RNI4EULD[28]  (.A(\counter[27]_net_1 ), .B(
        counter_c26), .C(\counter[28]_net_1 ), .Y(counter_c28));
    NOR2A un1_counter_2_0_I_19 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] ), .B(\counter[31]_net_1 )
        , .Y(\DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] ));
    OR2 \off_reg_RNI4UT6[6]  (.A(\off_reg[6]_net_1 ), .B(act_ctl_5_4), 
        .Y(\off_time[6] ));
    NOR2A un1_counter_0_I_46 (.A(\off_time[24] ), .B(
        \counter[24]_net_1 ), .Y(\ACT_LT3_E[0] ));
    NOR2A \off_reg_RNINR0Q[22]  (.A(\off_reg[22]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[22] ));
    GND GND_i (.Y(GND));
    DFN1C0 \counter[13]  (.D(counter_n13), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[13]_net_1 ));
    XNOR2 un1_counter_0_I_81 (.A(\counter[16]_net_1 ), .B(
        \off_time[16] ), .Y(\DWACT_BL_EQUAL_0_E_1[1] ));
    NOR2A un1_counter_0_I_90 (.A(\off_time[18] ), .B(
        \counter[18]_net_1 ), .Y(\ACT_LT4_E[5] ));
    XNOR2 un1_counter_0_I_74 (.A(\counter[11]_net_1 ), .B(
        \off_time[11] ), .Y(\DWACT_BL_EQUAL_0_E_2[1] ));
    NOR2B un1_counter_2_0_I_140 (.A(\DWACT_COMP0_E[2] ), .B(
        \DWACT_COMP0_E[1] ), .Y(I_140));
    OA1A un1_counter_0_I_36 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .C(N_43), .Y(N_47));
    XNOR2 un1_counter_0_I_66 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\DWACT_BL_EQUAL_0_E[8] ));
    AND3 un1_counter_0_I_17 (.A(\DWACT_BL_EQUAL_0_E_5[0] ), .B(
        \DWACT_BL_EQUAL_0_E_5[1] ), .C(\DWACT_BL_EQUAL_0_E_5[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] ));
    NOR3C \counter_RNI38793[5]  (.A(\counter[5]_net_1 ), .B(counter_c4)
        , .C(\counter[6]_net_1 ), .Y(counter_c6));
    DFN1E1C0 \off_reg[17]  (.D(off_div[17]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[17]_net_1 ));
    AX1C \counter_RNO_0[10]  (.A(\counter[9]_net_1 ), .B(counter_c8), 
        .C(\counter[10]_net_1 ), .Y(counter_n10_tz));
    DFN1C0 \counter[12]  (.D(counter_n12), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[12]_net_1 ));
    OR2A un1_counter_0_I_130 (.A(\off_time[4] ), .B(\counter[4]_net_1 )
        , .Y(N_5_0));
    NOR2B un1_counter_2_0_I_139 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E[2] )
        , .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ), .Y(
        \DWACT_COMP0_E[2] ));
    DFN1C0 \counter[27]  (.D(counter_n27), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[27]_net_1 ));
    OR2A un1_counter_0_I_96 (.A(\off_time[11] ), .B(
        \counter[11]_net_1 ), .Y(N_22));
    AOI1A un1_counter_0_I_49 (.A(\ACT_LT3_E[0] ), .B(\ACT_LT3_E[1] ), 
        .C(\ACT_LT3_E[2] ), .Y(\ACT_LT3_E[3] ));
    AX1C \counter_RNO_0[20]  (.A(\counter[19]_net_1 ), .B(counter_c18), 
        .C(\counter[20]_net_1 ), .Y(counter_n20_tz));
    DFN1C0 \counter[20]  (.D(counter_n20), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[20]_net_1 ));
    OA1A un1_counter_0_I_101 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .C(N_23), .Y(N_27));
    NOR3C \counter_RNI9T2D1[1]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .C(\counter[2]_net_1 ), .Y(counter_c2));
    NOR2A \off_reg_RNIMQ0Q[21]  (.A(\off_reg[21]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[21] ));
    DFN1E1C0 \off_reg[19]  (.D(off_div[19]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[19]_net_1 ));
    XNOR2 un1_counter_0_I_71 (.A(\counter[10]_net_1 ), .B(
        \off_time[10] ), .Y(\DWACT_BL_EQUAL_0_E_2[0] ));
    OR2A un1_counter_0_I_116 (.A(\off_time[6] ), .B(\counter[6]_net_1 )
        , .Y(N_12_0));
    AO1C un1_counter_0_I_39 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .C(N_45), .Y(N_50));
    XA1B \counter_RNO[17]  (.A(\counter[17]_net_1 ), .B(counter_c16), 
        .C(counter_N_3_0), .Y(counter_n17));
    XNOR2 un1_counter_0_I_69 (.A(\counter[16]_net_1 ), .B(
        \off_time[16] ), .Y(\DWACT_BL_EQUAL_0_E[6] ));
    XNOR2 un1_counter_0_I_112 (.A(\counter[9]_net_1 ), .B(
        \off_time[9] ), .Y(\DWACT_BL_EQUAL_0_E[4] ));
    OA1A un1_counter_0_I_105 (.A(N_26), .B(N_28), .C(N_27), .Y(N_31));
    DFN1C0 \counter[23]  (.D(counter_n23), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[23]_net_1 ));
    NOR2A \off_reg_RNILP0Q[20]  (.A(\off_reg[20]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[20] ));
    NOR2A \off_reg_RNI3TT6[5]  (.A(\off_reg[5]_net_1 ), .B(act_ctl_5_4)
        , .Y(\off_time[5] ));
    XA1B \counter_RNO[29]  (.A(\counter[29]_net_1 ), .B(counter_c28), 
        .C(counter_N_3_0), .Y(counter_n29));
    DFN1E1C0 \off_reg[25]  (.D(off_div[25]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[25]_net_1 ));
    NOR2B \counter_RNO_0[18]  (.A(counter_c16), .B(\counter[17]_net_1 )
        , .Y(counter_c17));
    DFN1C0 \counter[22]  (.D(counter_n22), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[22]_net_1 ));
    DFN1C0 \counter[15]  (.D(counter_n15), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[15]_net_1 ));
    AO1 un1_counter_0_I_107 (.A(\DWACT_CMPLE_PO0_DWACT_COMP0_E[1] ), 
        .B(\DWACT_CMPLE_PO0_DWACT_COMP0_E[2] ), .C(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] ));
    OR2A un1_counter_0_I_99 (.A(\off_time[14] ), .B(
        \counter[14]_net_1 ), .Y(N_25));
    AO1C un1_counter_2_0_I_122 (.A(\counter[7]_net_1 ), .B(I_20_0), .C(
        N_12), .Y(N_18));
    AND2 un1_counter_2_0_I_115 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] ));
    XNOR2 un1_counter_0_I_108 (.A(\counter[5]_net_1 ), .B(
        \off_time[5] ), .Y(\DWACT_BL_EQUAL_0_E_0[0] ));
    AX1C \counter_RNO_0[8]  (.A(\counter[7]_net_1 ), .B(counter_c6), 
        .C(\counter[8]_net_1 ), .Y(counter_n8_tz));
    AX1C \counter_RNO_0[28]  (.A(\counter[27]_net_1 ), .B(counter_c26), 
        .C(\counter[28]_net_1 ), .Y(counter_n28_tz));
    NOR2B \counter_RNI898M5[11]  (.A(counter_c10), .B(
        \counter[11]_net_1 ), .Y(counter_c11));
    VCC VCC_i (.Y(VCC));
    AO1C un1_counter_0_I_120 (.A(\off_time[6] ), .B(\counter[6]_net_1 )
        , .C(N_14_0), .Y(N_16_0));
    DFN1E1C0 \off_reg[31]  (.D(off_div[31]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[31]_net_1 ));
    NOR2A \counter_RNO_1[0]  (.A(primary_12_c), .B(\counter[0]_net_1 ), 
        .Y(counter_N_3_mux));
    XA1B \counter_RNO[14]  (.A(\counter[14]_net_1 ), .B(counter_c13), 
        .C(counter_N_3_0), .Y(counter_n14));
    NOR2B \counter_RNIAM467[14]  (.A(counter_c13), .B(
        \counter[14]_net_1 ), .Y(counter_c14));
    XNOR2 un1_counter_2_0_I_111 (.A(\counter[7]_net_1 ), .B(I_20_0), 
        .Y(\DWACT_BL_EQUAL_0_E[2] ));
    DFN1E1C0 \off_reg[7]  (.D(off_div[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[7]_net_1 ));
    NOR2B \counter_RNI1GULD[29]  (.A(counter_c28), .B(
        \counter[29]_net_1 ), .Y(counter_c29));
    DFN1C0 \counter[1]  (.D(\counter_RNO[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\counter[1]_net_1 ));
    XNOR2 un1_counter_0_I_2 (.A(\counter[19]_net_1 ), .B(
        \off_time[19] ), .Y(\DWACT_BL_EQUAL_0_E_5[0] ));
    NOR2A \counter_RNO[26]  (.A(counter_n26_tz), .B(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n26));
    NOR2A un1_counter_0_I_55 (.A(\off_time[19] ), .B(
        \counter[19]_net_1 ), .Y(N_34));
    AO1 un1_counter_0_I_139 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] ), .Y(\DWACT_COMP0_E_0[2] )
        );
    XA1B \counter_RNO[5]  (.A(\counter[5]_net_1 ), .B(counter_c4), .C(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n5));
    AO1C un1_counter_0_I_133 (.A(\counter[2]_net_1 ), .B(\off_time[2] )
        , .C(N_2), .Y(N_8_0));
    NOR2A un1_counter_2_0_I_132 (.A(N_3), .B(\counter[3]_net_1 ), .Y(
        N_7));
    OR2 \off_reg_RNI5VT6[7]  (.A(\off_reg[7]_net_1 ), .B(act_ctl_5_4), 
        .Y(\off_time[7] ));
    DFN1C0 \counter[25]  (.D(counter_n25), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[25]_net_1 ));
    AND2A un1_counter_0_I_87 (.A(\off_time[16] ), .B(
        \counter[16]_net_1 ), .Y(\ACT_LT4_E[2] ));
    XA1B \counter_RNO[3]  (.A(\counter[3]_net_1 ), .B(counter_c2), .C(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n3));
    DFN1E1C0 \off_reg[6]  (.D(off_div[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[6]_net_1 ));
    AND3 un1_counter_0_I_28 (.A(\DWACT_BL_EQUAL_0_E_4[0] ), .B(
        \DWACT_BL_EQUAL_0_E_4[1] ), .C(\DWACT_BL_EQUAL_0_E_4[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] ));
    NOR2A \off_reg_RNIRV0Q[26]  (.A(\off_reg[26]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[26] ));
    NOR2A \counter_RNO_0[0]  (.A(I_140_0), .B(\counter[0]_net_1 ), .Y(
        d_N_3_mux_4));
    OR2A un1_counter_0_I_50 (.A(\off_time[26] ), .B(
        \counter[26]_net_1 ), .Y(\ACT_LT3_E[4] ));
    DFN1C0 \counter[5]  (.D(counter_n5), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[5]_net_1 ));
    MX2A cur_pwm_RNO (.A(I_140_0), .B(I_140), .S(primary_12_c), .Y(
        cur_pwm_RNO_net_1));
    XNOR2 un1_counter_0_I_4 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(\DWACT_BL_EQUAL_0_E[10] ));
    XNOR2 un1_counter_0_I_23 (.A(\counter[27]_net_1 ), .B(
        \off_time[27] ), .Y(\DWACT_BL_EQUAL_0_E_4[0] ));
    NOR2A \counter_RNO[10]  (.A(counter_n10_tz), .B(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n10));
    AND3 un1_counter_0_I_77 (.A(\DWACT_BL_EQUAL_0_E_2[0] ), .B(
        \DWACT_BL_EQUAL_0_E_2[1] ), .C(\DWACT_BL_EQUAL_0_E_2[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] ));
    XNOR2 un1_counter_0_I_3 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .Y(\DWACT_BL_EQUAL_0_E[11] ));
    XA1B \counter_RNO[21]  (.A(\counter[21]_net_1 ), .B(counter_c20), 
        .C(counter_N_3_0), .Y(counter_n21));
    XNOR2 un1_counter_0_I_6 (.A(\counter[20]_net_1 ), .B(
        \off_time[20] ), .Y(\DWACT_BL_EQUAL_0_E_5[1] ));
    OR2A un1_counter_0_I_56 (.A(\off_time[23] ), .B(
        \counter[23]_net_1 ), .Y(N_35));
    AX1C \counter_RNO_0[24]  (.A(\counter[23]_net_1 ), .B(counter_c22), 
        .C(\counter[24]_net_1 ), .Y(counter_n24_tz));
    AND3 un1_counter_0_I_15 (.A(\DWACT_BL_EQUAL_0_E_0[6] ), .B(
        \DWACT_BL_EQUAL_0_E_0[7] ), .C(\DWACT_BL_EQUAL_0_E_0[8] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] ));
    NOR2B \counter_RNIRE268[16]  (.A(counter_c15), .B(
        \counter[16]_net_1 ), .Y(counter_c16));
    AND2A un1_counter_0_I_48 (.A(\off_time[25] ), .B(
        \counter[25]_net_1 ), .Y(\ACT_LT3_E[2] ));
    NOR2A un1_counter_0_I_129 (.A(\off_time[0] ), .B(
        \counter[0]_net_1 ), .Y(N_4));
    XNOR2 un1_counter_0_I_9 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(\DWACT_BL_EQUAL_0_E[12] ));
    AO1 un1_counter_0_I_140 (.A(\DWACT_COMP0_E_0[1] ), .B(
        \DWACT_COMP0_E_0[2] ), .C(\DWACT_COMP0_E[0] ), .Y(I_140_0));
    OR2A un1_counter_0_I_123 (.A(\counter[9]_net_1 ), .B(\off_time[9] )
        , .Y(N_19));
    DFN1C0 \counter[16]  (.D(counter_n16), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[16]_net_1 ));
    OR2A un1_counter_0_I_38 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(N_49));
    XA1B \counter_RNO[25]  (.A(\counter[25]_net_1 ), .B(counter_c24), 
        .C(counter_N_3_0), .Y(counter_n25));
    XNOR2 un1_counter_0_I_68 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\DWACT_BL_EQUAL_0_E[7] ));
    XNOR2 un1_act_ctl_I_14 (.A(N_4_0), .B(act_ctl_5_3), .Y(I_14_0));
    NOR2B \counter_RNO_0[31]  (.A(\counter[30]_net_1 ), .B(counter_c29)
        , .Y(\counter_RNO_0[31]_net_1 ));
    XNOR2 un1_counter_0_I_43 (.A(\counter[25]_net_1 ), .B(
        \off_time[25] ), .Y(\DWACT_BL_EQUAL_0_E_3[1] ));
    XOR2 un1_act_ctl_I_20 (.A(act_ctl_5_3), .B(N_2_0), .Y(I_20_0));
    AO1C un1_counter_0_I_59 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .C(N_32), .Y(N_38));
    DFN1E1C0 \off_reg[21]  (.D(off_div[21]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[21]_net_1 ));
    AO1C un1_counter_0_I_104 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .C(N_25), .Y(N_30));
    XNOR2 un1_counter_0_I_10 (.A(\counter[24]_net_1 ), .B(
        \off_time[24] ), .Y(\DWACT_BL_EQUAL_0_E_0[5] ));
    NOR2A \off_reg_RNISVVP[18]  (.A(\off_reg[18]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[18] ));
    NOR2A un1_counter_0_I_98 (.A(\off_time[10] ), .B(
        \counter[10]_net_1 ), .Y(N_24));
    NOR2A un1_counter_0_I_33 (.A(\off_time[27] ), .B(
        \counter[27]_net_1 ), .Y(N_44));
    OA1 un1_counter_0_I_63 (.A(N_41), .B(N_40), .C(N_39), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] ));
    NOR2A \counter_RNO[6]  (.A(counter_n6_tz), .B(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n6));
    XA1B \counter_RNO[30]  (.A(\counter[30]_net_1 ), .B(counter_c29), 
        .C(cur_pwm_RNIA74H44_0_net_1), .Y(counter_n30));
    MX2C cur_pwm_RNIA74H44 (.A(I_140_0), .B(I_140), .S(primary_12_c), 
        .Y(counter_N_3_0));
    XNOR2 un1_counter_0_I_110 (.A(\counter[8]_net_1 ), .B(
        \off_time[8] ), .Y(\DWACT_BL_EQUAL_0_E[3] ));
    DFN1E1C0 \off_reg[27]  (.D(off_div[27]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[27]_net_1 ));
    AND3 un1_counter_0_I_16 (.A(\DWACT_BL_EQUAL_0_E_3[3] ), .B(
        \DWACT_BL_EQUAL_0_E_2[4] ), .C(\DWACT_BL_EQUAL_0_E_0[5] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] ));
    NOR2A \off_reg_RNIQU0Q[25]  (.A(\off_reg[25]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[25] ));
    OR2A un1_counter_0_I_93 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\ACT_LT4_E[8] ));
    DFN1E1C0 \off_reg[8]  (.D(off_div[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[8]_net_1 ));
    DFN1C0 \counter[26]  (.D(counter_n26), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[26]_net_1 ));
    XA1B \counter_RNO[23]  (.A(\counter[23]_net_1 ), .B(counter_c22), 
        .C(counter_N_3_0), .Y(counter_n23));
    OA1 un1_counter_2_0_I_137 (.A(N_11), .B(N_10), .C(N_9), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] ));
    AO1C un1_counter_2_0_I_133 (.A(\counter[2]_net_1 ), .B(I_6), .C(
        \counter[1]_net_1 ), .Y(N_8));
    OR3A un1_act_ctl_I_19 (.A(act_ctl_5_0), .B(\DWACT_FDEC_E[2] ), .C(
        \DWACT_FDEC_E[0] ), .Y(N_2_0));
    DFN1C0 \counter[14]  (.D(counter_n14), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[14]_net_1 ));
    DFN1E1C0 \off_reg[29]  (.D(off_div[29]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[29]_net_1 ));
    AND3 un1_counter_2_0_I_18 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] ));
    DFN1E1C0 \off_reg[1]  (.D(off_div[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[1]_net_1 ));
    NOR2A \counter_RNO[22]  (.A(counter_n22_tz), .B(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n22));
    AO1C un1_counter_0_I_131 (.A(\off_time[1] ), .B(\counter[1]_net_1 )
        , .C(N_4), .Y(N_6_0));
    AND2 un1_counter_0_I_19 (.A(\DWACT_BL_EQUAL_0_E[12] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] ));
    XNOR2 un1_counter_0_I_42 (.A(\counter[26]_net_1 ), .B(
        \off_time[26] ), .Y(\DWACT_BL_EQUAL_0_E_3[2] ));
    AO1C un1_counter_0_I_135 (.A(\counter[3]_net_1 ), .B(\off_time[3] )
        , .C(N_5_0), .Y(N_10_0));
    DFN1E1C0 \off_reg[10]  (.D(off_div[10]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[10]_net_1 ));
    NOR2A un1_counter_0_I_85 (.A(\off_time[15] ), .B(
        \counter[15]_net_1 ), .Y(\ACT_LT4_E[0] ));
    DFN1C0 \counter[31]  (.D(counter_N_7), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[31]_net_1 ));
    NOR2A \off_reg_RNIRUVP[17]  (.A(\off_reg[17]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[17] ));
    OR2A un1_counter_0_I_32 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(N_43));
    OA1A un1_counter_0_I_62 (.A(N_36), .B(N_38), .C(N_37), .Y(N_41));
    OR3A un1_act_ctl_I_13 (.A(act_ctl_5_0), .B(act_ctl_5_0), .C(
        \DWACT_FDEC_E[0] ), .Y(N_4_0));
    OA1 un1_counter_0_I_137 (.A(N_11_0), .B(N_10_0), .C(N_9_0), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] ));
    AO1 un1_counter_0_I_138 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] ));
    NOR2A un1_counter_0_I_92 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\ACT_LT4_E[7] ));
    DFN1C0 \counter[24]  (.D(counter_n24), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[24]_net_1 ));
    OR2A un1_counter_0_I_119 (.A(\off_time[9] ), .B(\counter[9]_net_1 )
        , .Y(N_15));
    NOR3 un1_counter_2_0_I_14 (.A(\counter[29]_net_1 ), .B(
        \counter[30]_net_1 ), .C(\counter[28]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] ));
    MX2C cur_pwm_RNIA74H44_0 (.A(I_140_0), .B(I_140), .S(primary_12_c), 
        .Y(cur_pwm_RNIA74H44_0_net_1));
    AND3 un1_counter_2_0_I_78 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ));
    XNOR2 un1_counter_0_I_80 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\DWACT_BL_EQUAL_0_E_1[2] ));
    XNOR2 un1_counter_0_I_5 (.A(\counter[27]_net_1 ), .B(
        \off_time[27] ), .Y(\DWACT_BL_EQUAL_0_E_0[8] ));
    AND3 un1_counter_0_I_113 (.A(\DWACT_BL_EQUAL_0_E_0[0] ), .B(
        \DWACT_BL_EQUAL_0_E_0[1] ), .C(\DWACT_BL_EQUAL_0_E_0[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] ));
    XNOR2 un1_counter_0_I_24 (.A(\counter[28]_net_1 ), .B(
        \off_time[28] ), .Y(\DWACT_BL_EQUAL_0_E_4[1] ));
    NOR2A \counter_RNO[4]  (.A(counter_n4_tz), .B(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n4));
    AND3 un1_counter_0_I_75 (.A(\DWACT_BL_EQUAL_0_E[6] ), .B(
        \DWACT_BL_EQUAL_0_E[7] ), .C(\DWACT_BL_EQUAL_0_E[8] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] ));
    DFN1E1C0 \off_reg[14]  (.D(off_div[14]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[14]_net_1 ));
    NOR2A \off_reg_RNIUNT6[0]  (.A(\off_reg[0]_net_1 ), .B(act_ctl_5_4)
        , .Y(\off_time[0] ));
    AO1C un1_counter_2_0_I_120 (.A(I_17_0), .B(\counter[6]_net_1 ), .C(
        N_14), .Y(N_16));
    XA1B \counter_RNO[18]  (.A(\counter[18]_net_1 ), .B(counter_c17), 
        .C(counter_N_3_0), .Y(counter_n18));
    NOR3C \counter_RNIBOU5B[22]  (.A(\counter[21]_net_1 ), .B(
        counter_c20), .C(\counter[22]_net_1 ), .Y(counter_c22));
    NOR3 un1_counter_2_0_I_15 (.A(\counter[26]_net_1 ), .B(
        \counter[27]_net_1 ), .C(\counter[25]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] ));
    OR2A un1_counter_0_I_86 (.A(\off_time[16] ), .B(
        \counter[16]_net_1 ), .Y(\ACT_LT4_E[1] ));
    OA1A un1_counter_0_I_58 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .C(N_33), .Y(N_37));
    OA1A un1_counter_0_I_121 (.A(\counter[8]_net_1 ), .B(\off_time[8] )
        , .C(N_13_0), .Y(N_17_0));
    OR2 \off_reg_RNI2ST6[4]  (.A(\off_reg[4]_net_1 ), .B(act_ctl_5_4), 
        .Y(\off_time[4] ));
    AND2 un1_counter_2_0_I_20 (.A(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] ), .B(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] ), .Y(
        \DWACT_COMP0_E[1] ));
    AX1C \counter_RNO_0[26]  (.A(\counter[25]_net_1 ), .B(counter_c24), 
        .C(\counter[26]_net_1 ), .Y(counter_n26_tz));
    XA1B \counter_RNO[27]  (.A(\counter[27]_net_1 ), .B(counter_c26), 
        .C(counter_N_3_0), .Y(counter_n27));
    OA1A un1_counter_0_I_125 (.A(N_16_0), .B(N_18_0), .C(N_17_0), .Y(
        N_21_0));
    AX1C \counter_RNO_0[6]  (.A(\counter[5]_net_1 ), .B(counter_c4), 
        .C(\counter[6]_net_1 ), .Y(counter_n6_tz));
    XNOR2 un1_counter_0_I_70 (.A(\counter[15]_net_1 ), .B(
        \off_time[15] ), .Y(\DWACT_BL_EQUAL_0_E[5] ));
    OA1 un1_counter_0_I_106 (.A(N_31), .B(N_30), .C(N_29), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] ));
    NOR3C \counter_RNI04V5A[19]  (.A(\counter[19]_net_1 ), .B(
        counter_c18), .C(\counter[20]_net_1 ), .Y(counter_c20));
    OR2A un1_act_ctl_I_15 (.A(act_ctl_5_3), .B(act_ctl_5_3), .Y(
        \DWACT_FDEC_E[1] ));
    DFN1E1C0 \off_reg[18]  (.D(off_div[18]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[18]_net_1 ));
    AO1C un1_counter_0_I_102 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .C(N_22), .Y(N_28));
    OR2A un1_counter_2_0_I_117 (.A(\counter[7]_net_1 ), .B(I_20_0), .Y(
        N_13));
    AND3 un1_counter_2_0_I_113 (.A(\DWACT_BL_EQUAL_0_E[0] ), .B(
        \DWACT_BL_EQUAL_0_E[1] ), .C(\DWACT_BL_EQUAL_0_E[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ));
    XNOR2 un1_counter_0_I_44 (.A(\counter[24]_net_1 ), .B(
        \off_time[24] ), .Y(\DWACT_BL_EQUAL_0_E_3[0] ));
    OR2A un1_counter_0_I_53 (.A(\off_time[20] ), .B(
        \counter[20]_net_1 ), .Y(N_32));
    NOR2A \off_reg_RNI60U6[8]  (.A(\off_reg[8]_net_1 ), .B(act_ctl_5_4)
        , .Y(\off_time[8] ));
    OR2A un1_counter_0_I_127 (.A(\off_time[1] ), .B(\counter[1]_net_1 )
        , .Y(N_2));
    XOR2 un1_act_ctl_I_17 (.A(act_ctl_5_3), .B(N_3_1), .Y(I_17_0));
    NOR2A \off_reg_RNI71U6[9]  (.A(\off_reg[9]_net_1 ), .B(act_ctl_5_4)
        , .Y(\off_time[9] ));
    XNOR2 un1_act_ctl_I_12 (.A(N_5), .B(act_ctl_5_3), .Y(I_12_0));
    NOR2A un1_counter_2_0_I_130 (.A(I_12_0), .B(\counter[4]_net_1 ), 
        .Y(N_10));
    OR2A un1_counter_0_I_34 (.A(\off_time[31] ), .B(
        \counter[31]_net_1 ), .Y(N_45));
    OR2A un1_counter_0_I_128 (.A(\counter[2]_net_1 ), .B(\off_time[2] )
        , .Y(N_3_0));
    OR2A un1_counter_0_I_89 (.A(\off_time[17] ), .B(
        \counter[17]_net_1 ), .Y(\ACT_LT4_E[4] ));
    AO1 un1_counter_0_I_64 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] ));
    DFN1E1C0 \off_reg[16]  (.D(off_div[16]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[16]_net_1 ));
    AND3 un1_counter_0_I_76 (.A(\DWACT_BL_EQUAL_0_E_1[3] ), .B(
        \DWACT_BL_EQUAL_0_E_0[4] ), .C(\DWACT_BL_EQUAL_0_E[5] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] ));
    XNOR2 un1_counter_0_I_1 (.A(\counter[23]_net_1 ), .B(
        \off_time[23] ), .Y(\DWACT_BL_EQUAL_0_E_2[4] ));
    OR2A un1_counter_2_0_I_134 (.A(\counter[4]_net_1 ), .B(I_12_0), .Y(
        N_9));
    DFN1E1C0 \off_reg[30]  (.D(off_div[30]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[30]_net_1 ));
    NOR3 un1_counter_2_0_I_75 (.A(\counter[17]_net_1 ), .B(
        \counter[18]_net_1 ), .C(\counter[16]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] ));
    NOR2A \counter_RNO[24]  (.A(counter_n24_tz), .B(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n24));
    DFN1C0 \counter[7]  (.D(counter_n7), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[7]_net_1 ));
    AOI1A un1_counter_0_I_94 (.A(\ACT_LT4_E[7] ), .B(\ACT_LT4_E[8] ), 
        .C(\ACT_LT4_E[5] ), .Y(\ACT_LT4_E[10] ));
    DFN1C0 \counter[30]  (.D(counter_n30), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[30]_net_1 ));
    NOR3C \counter_RNI5GSF1[10]  (.A(\counter[15]_net_1 ), .B(
        \counter[10]_net_1 ), .C(\counter[17]_net_1 ), .Y(
        counter_m6_0_a2_4));
    OA1 un1_counter_0_I_41 (.A(N_51), .B(N_50), .C(N_49), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] ));
    OR3 un1_act_ctl_I_16 (.A(\DWACT_FDEC_E[0] ), .B(\DWACT_FDEC_E[1] ), 
        .C(act_ctl_5_0), .Y(N_3_1));
    AND3 un1_counter_0_I_18 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] ));
    NOR2B \counter_RNIDKTV[13]  (.A(\counter[13]_net_1 ), .B(
        \counter[14]_net_1 ), .Y(counter_m6_0_a2_2));
    OR2A un1_counter_0_I_31 (.A(\off_time[28] ), .B(
        \counter[28]_net_1 ), .Y(N_42));
    XNOR2 un1_counter_2_0_I_108 (.A(\counter[5]_net_1 ), .B(I_14_0), 
        .Y(\DWACT_BL_EQUAL_0_E[0] ));
    AO1C un1_counter_0_I_61 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .C(N_35), .Y(N_40));
    MX2 \counter_RNO[0]  (.A(d_N_3_mux_4), .B(I_140), .S(
        counter_N_3_mux), .Y(\counter_RNO[0]_net_1 ));
    XNOR2 un1_counter_0_I_79 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\DWACT_BL_EQUAL_0_E_0[3] ));
    NOR2A \off_reg_RNIORVP[14]  (.A(\off_reg[14]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[14] ));
    NOR3C \counter_RNIKH965[10]  (.A(\counter[9]_net_1 ), .B(
        counter_c8), .C(\counter[10]_net_1 ), .Y(counter_c10));
    DFN1E1C0 \off_reg[3]  (.D(off_div[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[3]_net_1 ));
    DFN1E1C0 \off_reg[0]  (.D(off_div[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[0]_net_1 ));
    NOR3C \counter_RNIK05B2[3]  (.A(\counter[3]_net_1 ), .B(counter_c2)
        , .C(\counter[4]_net_1 ), .Y(counter_c4));
    OR3 un1_act_ctl_I_18 (.A(act_ctl_5_i), .B(act_ctl_5_0), .C(
        act_ctl_5_0), .Y(\DWACT_FDEC_E[2] ));
    NOR2A \off_reg_RNIQTVP[16]  (.A(\off_reg[16]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[16] ));
    NOR2B \counter_RNIT1766[12]  (.A(counter_c11), .B(
        \counter[12]_net_1 ), .Y(counter_c12));
    NOR2A un1_counter_2_0_I_126 (.A(N_21), .B(\counter[9]_net_1 ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ));
    OR2A un1_counter_0_I_134 (.A(\counter[4]_net_1 ), .B(\off_time[4] )
        , .Y(N_9_0));
    XNOR2 un1_counter_0_I_13 (.A(\counter[28]_net_1 ), .B(
        \off_time[28] ), .Y(\DWACT_BL_EQUAL_0_E[9] ));
    NOR2A \off_reg_RNIPSVP[15]  (.A(\off_reg[15]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[15] ));
    OR2 \off_reg_RNI1RT6[3]  (.A(\off_reg[3]_net_1 ), .B(act_ctl_5_4), 
        .Y(\off_time[3] ));
    NOR2A un1_counter_0_I_91 (.A(\ACT_LT4_E[4] ), .B(\ACT_LT4_E[5] ), 
        .Y(\ACT_LT4_E[6] ));
    AOI1A un1_counter_0_I_52 (.A(\ACT_LT3_E[3] ), .B(\ACT_LT3_E[4] ), 
        .C(\ACT_LT3_E[5] ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] ));
    NOR2A \counter_RNO_2[1]  (.A(primary_12_c), .B(I_140), .Y(
        counter_N_7_0));
    NOR2A \counter_RNO[20]  (.A(counter_n20_tz), .B(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n20));
    NOR3C \counter_RNIQGU5C[24]  (.A(\counter[23]_net_1 ), .B(
        counter_c22), .C(\counter[24]_net_1 ), .Y(counter_c24));
    NOR3C \counter_RNIGB069[9]  (.A(\counter[9]_net_1 ), .B(counter_c8)
        , .C(counter_m6_0_a2_7), .Y(counter_c18));
    DFN1E1C0 \off_reg[13]  (.D(off_div[13]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[13]_net_1 ));
    OR2A un1_counter_2_0_I_128 (.A(\counter[2]_net_1 ), .B(I_6), .Y(
        N_3));
    XNOR2 un1_counter_0_I_27 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(\DWACT_BL_EQUAL_0_E_1[4] ));
    XNOR2 un1_counter_0_I_111 (.A(\counter[7]_net_1 ), .B(
        \off_time[7] ), .Y(\DWACT_BL_EQUAL_0_E_0[2] ));
    OA1A un1_counter_2_0_I_136 (.A(N_6), .B(N_8), .C(N_7), .Y(N_11));
    NOR2B \counter_RNI9GTV[11]  (.A(\counter[11]_net_1 ), .B(
        \counter[12]_net_1 ), .Y(counter_m6_0_a2_1));
    AND2 un1_counter_0_I_115 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] ));
    DFN1E1C0 \off_reg[4]  (.D(off_div[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[4]_net_1 ));
    XNOR2 un1_counter_0_I_8 (.A(\counter[25]_net_1 ), .B(
        \off_time[25] ), .Y(\DWACT_BL_EQUAL_0_E_0[6] ));
    DFN1E1C0 \off_reg[20]  (.D(off_div[20]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[20]_net_1 ));
    NOR2A \counter_RNO[2]  (.A(counter_n2_tz), .B(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n2));
    DFN1C0 \counter[9]  (.D(counter_n9), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[9]_net_1 ));
    NOR3 un1_counter_2_0_I_16 (.A(\counter[24]_net_1 ), .B(
        \counter[23]_net_1 ), .C(\counter[22]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] ));
    NOR2 un1_counter_2_0_I_114 (.A(\counter[8]_net_1 ), .B(
        \counter[9]_net_1 ), .Y(\DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ));
    OR2A un1_counter_0_I_117 (.A(\counter[7]_net_1 ), .B(\off_time[7] )
        , .Y(N_13_0));
    XA1B \counter_RNO[19]  (.A(\counter[19]_net_1 ), .B(counter_c18), 
        .C(counter_N_3_0), .Y(counter_n19));
    AO1C un1_counter_0_I_124 (.A(\counter[8]_net_1 ), .B(\off_time[8] )
        , .C(N_15), .Y(N_20));
    NOR2A un1_counter_0_I_118 (.A(\off_time[5] ), .B(
        \counter[5]_net_1 ), .Y(N_14_0));
    XNOR2 un1_counter_0_I_12 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .Y(\DWACT_BL_EQUAL_0_E_5[2] ));
    AO1 un1_counter_2_0_I_138 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] )
        , .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] ));
    XA1B \counter_RNO[9]  (.A(\counter[9]_net_1 ), .B(counter_c8), .C(
        cur_pwm_RNIA74H44_0_net_1), .Y(counter_n9));
    DFN1E1C0 \off_reg[12]  (.D(off_div[12]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[12]_net_1 ));
    AOI1A un1_counter_0_I_88 (.A(\ACT_LT4_E[0] ), .B(\ACT_LT4_E[1] ), 
        .C(\ACT_LT4_E[2] ), .Y(\ACT_LT4_E[3] ));
    OR2A un1_counter_0_I_47 (.A(\off_time[25] ), .B(
        \counter[25]_net_1 ), .Y(\ACT_LT3_E[1] ));
    DFN1C0 \counter[8]  (.D(counter_n8), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[8]_net_1 ));
    NOR2A \off_reg_RNIVUFT[31]  (.A(\off_reg[31]_net_1 ), .B(act_ctl_5)
        , .Y(\off_time[31] ));
    OR2A un1_counter_0_I_54 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .Y(N_33));
    AO1C un1_counter_0_I_37 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .C(N_42), .Y(N_48));
    XNOR2 un1_counter_0_I_7 (.A(\counter[26]_net_1 ), .B(
        \off_time[26] ), .Y(\DWACT_BL_EQUAL_0_E_0[7] ));
    XNOR2 un1_counter_0_I_67 (.A(\counter[14]_net_1 ), .B(
        \off_time[14] ), .Y(\DWACT_BL_EQUAL_0_E_0[4] ));
    DFN1C0 \counter[18]  (.D(counter_n18), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[18]_net_1 ));
    AO1C un1_counter_0_I_100 (.A(\off_time[11] ), .B(
        \counter[11]_net_1 ), .C(N_24), .Y(N_26));
    DFN1E1C0 \off_reg[24]  (.D(off_div[24]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[24]_net_1 ));
    AND3 un1_counter_0_I_83 (.A(\DWACT_BL_EQUAL_0_E_1[0] ), .B(
        \DWACT_BL_EQUAL_0_E_1[1] ), .C(\DWACT_BL_EQUAL_0_E_1[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] ));
    XA1B \counter_RNO[16]  (.A(\counter[16]_net_1 ), .B(counter_c15), 
        .C(counter_N_3_0), .Y(counter_n16));
    DFN1C0 \counter[0]  (.D(\counter_RNO[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\counter[0]_net_1 ));
    NOR3 un1_counter_2_0_I_76 (.A(\counter[15]_net_1 ), .B(
        \counter[14]_net_1 ), .C(\counter[13]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] ));
    OR2A un1_counter_0_I_97 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .Y(N_23));
    NOR2A \off_reg_RNIOS0Q[23]  (.A(\off_reg[23]_net_1 ), .B(
        act_ctl_5_9), .Y(\off_time[23] ));
    
endmodule


module spi_clk_11s_0(
       cur_clk,
       n_rst_c,
       clk_c
    );
output cur_clk;
input  n_rst_c;
input  clk_c;

    wire N_8, \counter[1]_net_1 , \counter[0]_net_1 , N_6, 
        \counter[3]_net_1 , \DWACT_FINC_E[0] , cur_clk5_5, cur_clk5_3, 
        \counter[6]_net_1 , cur_clk5_4, cur_clk5_1, \counter[7]_net_1 , 
        \counter[8]_net_1 , \counter[4]_net_1 , \counter[5]_net_1 , 
        \counter[2]_net_1 , cur_clk_RNO_net_1, \counter_3[1] , I_5, 
        \counter_3[0] , \counter_3[3] , I_9, I_7, I_12, I_14, I_17, 
        I_20, I_23, N_2, \DWACT_FINC_E[2] , \DWACT_FINC_E[3] , N_3, 
        N_4, \DWACT_FINC_E[1] , N_5, N_7, GND, VCC;
    
    NOR2B un3_counter_I_6 (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(N_8));
    AND3 un3_counter_I_19 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\counter[6]_net_1 ), .Y(N_3));
    XOR2 un3_counter_I_20 (.A(N_3), .B(\counter[7]_net_1 ), .Y(I_20));
    NOR3A \counter_RNIQNI8[8]  (.A(cur_clk5_1), .B(\counter[7]_net_1 ), 
        .C(\counter[8]_net_1 ), .Y(cur_clk5_4));
    DFN1C0 \counter[2]  (.D(I_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[2]_net_1 ));
    NOR2A \counter_RNIP794[4]  (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(cur_clk5_3));
    DFN1C0 \counter[7]  (.D(I_20), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[7]_net_1 ));
    AND3 un3_counter_I_13 (.A(\DWACT_FINC_E[0] ), .B(
        \counter[3]_net_1 ), .C(\counter[4]_net_1 ), .Y(N_5));
    AOI1 \counter_RNO[0]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(
        \counter[0]_net_1 ), .Y(\counter_3[0] ));
    DFN1C0 \counter[6]  (.D(I_17), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[6]_net_1 ));
    VCC VCC_i (.Y(VCC));
    XOR2 un3_counter_I_12 (.A(N_6), .B(\counter[4]_net_1 ), .Y(I_12));
    DFN1C0 \counter[8]  (.D(I_23), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[8]_net_1 ));
    XOR2 un3_counter_I_23 (.A(N_2), .B(\counter[8]_net_1 ), .Y(I_23));
    AOI1B \counter_RNO[1]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(I_5), 
        .Y(\counter_3[1] ));
    AND3 un3_counter_I_22 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\DWACT_FINC_E[3] ), .Y(N_2));
    XOR2 un3_counter_I_7 (.A(N_8), .B(\counter[2]_net_1 ), .Y(I_7));
    NOR2B un3_counter_I_11 (.A(\counter[3]_net_1 ), .B(
        \DWACT_FINC_E[0] ), .Y(N_6));
    AND3 un3_counter_I_16 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[1] )
        , .C(\counter[5]_net_1 ), .Y(N_4));
    DFN1C0 \counter[4]  (.D(I_12), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[4]_net_1 ));
    XOR2 un3_counter_I_17 (.A(N_4), .B(\counter[6]_net_1 ), .Y(I_17));
    NOR2 \counter_RNIP794[2]  (.A(\counter[5]_net_1 ), .B(
        \counter[2]_net_1 ), .Y(cur_clk5_1));
    DFN1C0 \counter[5]  (.D(I_14), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[5]_net_1 ));
    AND3 un3_counter_I_8 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(N_7));
    GND GND_i (.Y(GND));
    AX1C cur_clk_RNO (.A(cur_clk5_4), .B(cur_clk5_5), .C(cur_clk), .Y(
        cur_clk_RNO_net_1));
    AOI1B \counter_RNO[3]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(I_9), 
        .Y(\counter_3[3] ));
    AND2 un3_counter_I_21 (.A(\counter[6]_net_1 ), .B(
        \counter[7]_net_1 ), .Y(\DWACT_FINC_E[3] ));
    DFN1C0 \counter[1]  (.D(\counter_3[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[1]_net_1 ));
    DFN1C0 \counter[3]  (.D(\counter_3[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[3]_net_1 ));
    NOR3B \counter_RNIIFI8[6]  (.A(\counter[1]_net_1 ), .B(cur_clk5_3), 
        .C(\counter[6]_net_1 ), .Y(cur_clk5_5));
    AND2 un3_counter_I_15 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(\DWACT_FINC_E[1] ));
    XOR2 un3_counter_I_9 (.A(N_7), .B(\counter[3]_net_1 ), .Y(I_9));
    DFN1C0 cur_clk_inst_1 (.D(cur_clk_RNO_net_1), .CLK(clk_c), .CLR(
        n_rst_c), .Q(cur_clk));
    XOR2 un3_counter_I_14 (.A(N_5), .B(\counter[5]_net_1 ), .Y(I_14));
    XOR2 un3_counter_I_5 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .Y(I_5));
    AND3 un3_counter_I_10 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(
        \DWACT_FINC_E[0] ));
    DFN1C0 \counter[0]  (.D(\counter_3[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[0]_net_1 ));
    AND3 un3_counter_I_18 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .C(\counter[5]_net_1 ), .Y(
        \DWACT_FINC_E[2] ));
    
endmodule


module PID_controller_Z2(
       choose_0_0,
       choose,
       LED_15,
       LED_c,
       LED_5,
       LED_FB,
       LED_33,
       LED_12,
       primary_12_c,
       act_ctl_5_7,
       act_ctl_5_3,
       act_ctl_5_4,
       act_ctl_5_9,
       act_ctl_5,
       act_ctl_5_8,
       act_ctl_5_0,
       act_ctl_5_i,
       din_12_c,
       cs_i_1_i,
       cur_clk,
       clk_c,
       n_rst_c
    );
input  choose_0_0;
input  [2:0] choose;
input  [7:6] LED_15;
output [7:6] LED_c;
input  [7:6] LED_5;
input  [7:6] LED_FB;
input  [7:6] LED_33;
output [5:0] LED_12;
output primary_12_c;
input  act_ctl_5_7;
input  act_ctl_5_3;
input  act_ctl_5_4;
input  act_ctl_5_9;
input  act_ctl_5;
input  act_ctl_5_8;
input  act_ctl_5_0;
input  act_ctl_5_i;
input  din_12_c;
output cs_i_1_i;
output cur_clk;
input  clk_c;
input  n_rst_c;

    wire \state[1] , \state[0] , pwm_chg, sig_prev, sig_old_i_0, 
        N_46_1, avg_done, sig_old_i_0_0, sig_prev_0, sum_rdy, 
        deriv_enable, calc_avg, calc_int, pwm_enable, sum_enable, 
        calc_error, avg_enable, int_enable, pwm_chg_0, avg_enable_0, 
        avg_enable_1, \cur_vd[0] , \cur_vd[1] , \cur_vd[2] , 
        \cur_vd[3] , \cur_vd[4] , \cur_vd[5] , \cur_vd[6] , 
        \cur_vd[7] , \cur_vd[8] , \cur_vd[9] , \cur_vd[10] , 
        \cur_vd[11] , \avg_new[0] , \avg_new[1] , \avg_new[2] , 
        \avg_new[3] , \avg_new[4] , \avg_new[5] , \avg_new[6] , 
        \avg_new[7] , \avg_new[8] , \avg_new[9] , \avg_new[10] , 
        \avg_new[11] , \avg_old[0] , \avg_old[1] , \avg_old[2] , 
        \avg_old[3] , \avg_old[4] , \avg_old[5] , \avg_old[6] , 
        \avg_old[7] , \avg_old[8] , \avg_old[9] , \avg_old[10] , 
        \avg_old[11] , \cur_error[0] , \cur_error[1] , \cur_error[2] , 
        \cur_error[3] , \cur_error[4] , \cur_error[5] , \cur_error[6] , 
        \cur_error[7] , \cur_error[8] , \cur_error[9] , 
        \cur_error[10] , \cur_error[11] , \cur_error[12] , 
        \LED_12_i[5] , \LED_12[6] , \LED_12[7] , \average[2] , 
        \average[3] , \average[4] , \average[5] , \average[6] , 
        \sr_old[0] , \sr_old[1] , \sr_old[2] , \sr_old[3] , 
        \sr_old[4] , \sr_old[5] , \sr_old[6] , \sr_old[7] , 
        \sr_old[8] , \sr_old[9] , \sr_old[10] , \sr_old[11] , 
        \sr_old[12] , \sr_new[0] , \sr_new[1] , \sr_new[2] , 
        \sr_new[3] , \sr_new[4] , \sr_new[5] , \sr_new[6] , 
        \sr_new[7] , \sr_new[8] , \sr_new[9] , \sr_new[10] , 
        \sr_new[11] , \sr_new[12] , \sr_prev[0] , \sr_prev[1] , 
        \sr_prev[2] , \sr_prev[3] , \sr_prev[4] , \sr_prev[5] , 
        \sr_prev[6] , \sr_prev[7] , \sr_prev[8] , \sr_prev[9] , 
        \sr_prev[10] , \sr_prev[11] , \sr_prev[12] , \sr_new_0[12] , 
        \sr_new_1[12] , \integral[6] , \integral[7] , \integral[8] , 
        \integral[9] , \integral[10] , \integral[11] , \integral[12] , 
        \integral[13] , \integral[14] , \integral[15] , \integral[16] , 
        \integral[17] , \integral[18] , \integral[19] , \integral[20] , 
        \integral[21] , \integral[22] , \integral[23] , \integral[24] , 
        \integral[25] , \integral_i[24] , \integral_i[25] , 
        \integral_0[25] , \integral_1[25] , \derivative[12] , 
        \sum[39] , \sum[14] , \sum[19] , \sum[20] , \sum[22] , 
        \sum[13] , \sum[18] , \sum[17] , \sum[23] , \sum[21] , 
        \sum[16] , \sum[15] , \sum[12] , \sum[11] , \sum[6] , 
        \sum[10] , \sum[9] , \sum[5] , \sum[8] , \sum[7] , \sum[4] , 
        \sum[2] , \sum[1] , \sum[0] , \sum[3] , \sum_0[39] , 
        \sum_1[39] , \sum_2[39] , vd_done, \off_div[0] , \off_div[1] , 
        \off_div[2] , \off_div[3] , \off_div[4] , \off_div[5] , 
        \off_div[6] , \off_div[7] , \off_div[8] , \off_div[9] , 
        \off_div[10] , \off_div[11] , \off_div[12] , \off_div[13] , 
        \off_div[14] , \off_div[15] , \off_div[16] , \off_div[17] , 
        \off_div[18] , \off_div[19] , \off_div[20] , \off_div[21] , 
        \off_div[22] , \off_div[23] , \off_div[24] , \off_div[25] , 
        \off_div[26] , \off_div[27] , \off_div[28] , \off_div[29] , 
        \off_div[30] , \off_div[31] , GND, VCC;
    
    pwm_ctl_200s_32s_13s_0_1_2_1 PWM_CTL (.sum_8(\sum[8] ), .sum_39(
        \sum[39] ), .sum_12(\sum[12] ), .sum_14(\sum[14] ), .sum_15(
        \sum[15] ), .sum_16(\sum[16] ), .sum_17(\sum[17] ), .sum_18(
        \sum[18] ), .sum_21(\sum[21] ), .sum_22(\sum[22] ), .sum_23(
        \sum[23] ), .sum_9(\sum[9] ), .sum_10(\sum[10] ), .sum_19(
        \sum[19] ), .sum_11(\sum[11] ), .sum_20(\sum[20] ), .sum_13(
        \sum[13] ), .sum_1_d0(\sum[1] ), .sum_0_d0(\sum[0] ), 
        .sum_2_d0(\sum[2] ), .sum_7(\sum[7] ), .sum_6(\sum[6] ), 
        .sum_3(\sum[3] ), .sum_5(\sum[5] ), .sum_4(\sum[4] ), .sum_0_0(
        \sum_0[39] ), .off_div({\off_div[31] , \off_div[30] , 
        \off_div[29] , \off_div[28] , \off_div[27] , \off_div[26] , 
        \off_div[25] , \off_div[24] , \off_div[23] , \off_div[22] , 
        \off_div[21] , \off_div[20] , \off_div[19] , \off_div[18] , 
        \off_div[17] , \off_div[16] , \off_div[15] , \off_div[14] , 
        \off_div[13] , \off_div[12] , \off_div[11] , \off_div[10] , 
        \off_div[9] , \off_div[8] , \off_div[7] , \off_div[6] , 
        \off_div[5] , \off_div[4] , \off_div[3] , \off_div[2] , 
        \off_div[1] , \off_div[0] }), .sum_1_0(\sum_1[39] ), .sum_2_0(
        \sum_2[39] ), .state({\state[1] , \state[0] }), .n_rst_c(
        n_rst_c), .clk_c(clk_c), .pwm_enable(pwm_enable));
    integral_calc_13s_4 AVG_CALC (.avg_old({\avg_old[11] , 
        \avg_old[10] , \avg_old[9] , \avg_old[8] , \avg_old[7] , 
        \avg_old[6] , \avg_old[5] , \avg_old[4] , \avg_old[3] , 
        \avg_old[2] , \avg_old[1] , \avg_old[0] }), .avg_new({
        \avg_new[11] , \avg_new[10] , \avg_new[9] , \avg_new[8] , 
        \avg_new[7] , \avg_new[6] , \avg_new[5] , \avg_new[4] , 
        \avg_new[3] , \avg_new[2] , \avg_new[1] , \avg_new[0] }), 
        .LED_33({LED_33[7], LED_33[6]}), .LED_FB({LED_FB[7], LED_FB[6]})
        , .LED_5({LED_5[7], LED_5[6]}), .LED_c({LED_c[7], LED_c[6]}), 
        .LED_15({LED_15[7], LED_15[6]}), .choose({choose[2], choose[1], 
        choose[0]}), .choose_0_0(choose_0_0), .LED_12({\LED_12[7] , 
        \LED_12[6] , LED_12[5], LED_12[4], LED_12[3], LED_12[2], 
        LED_12[1], LED_12[0]}), .average({\average[6] , \average[5] , 
        \average[4] , \average[3] , \average[2] }), .LED_12_i_0(
        \LED_12_i[5] ), .avg_done(avg_done), .calc_avg(calc_avg), 
        .n_rst_c(n_rst_c), .clk_c(clk_c));
    error_sr_13s_5s AVGSR (.cur_vd({\cur_vd[11] , \cur_vd[10] , 
        \cur_vd[9] , \cur_vd[8] , \cur_vd[7] , \cur_vd[6] , 
        \cur_vd[5] , \cur_vd[4] , \cur_vd[3] , \cur_vd[2] , 
        \cur_vd[1] , \cur_vd[0] }), .avg_new({\avg_new[11] , 
        \avg_new[10] , \avg_new[9] , \avg_new[8] , \avg_new[7] , 
        \avg_new[6] , \avg_new[5] , \avg_new[4] , \avg_new[3] , 
        \avg_new[2] , \avg_new[1] , \avg_new[0] }), .avg_old({
        \avg_old[11] , \avg_old[10] , \avg_old[9] , \avg_old[8] , 
        \avg_old[7] , \avg_old[6] , \avg_old[5] , \avg_old[4] , 
        \avg_old[3] , \avg_old[2] , \avg_old[1] , \avg_old[0] }), 
        .avg_enable_1(avg_enable_1), .avg_enable_0(avg_enable_0), 
        .avg_enable(avg_enable), .n_rst_c(n_rst_c), .clk_c(clk_c));
    error_sr_13s_64s INTSR (.sr_old({\sr_old[12] , \sr_old[11] , 
        \sr_old[10] , \sr_old[9] , \sr_old[8] , \sr_old[7] , 
        \sr_old[6] , \sr_old[5] , \sr_old[4] , \sr_old[3] , 
        \sr_old[2] , \sr_old[1] , \sr_old[0] }), .sr_new({\sr_new[12] , 
        \sr_new[11] , \sr_new[10] , \sr_new[9] , \sr_new[8] , 
        \sr_new[7] , \sr_new[6] , \sr_new[5] , \sr_new[4] , 
        \sr_new[3] , \sr_new[2] , \sr_new[1] , \sr_new[0] }), 
        .cur_error({\cur_error[12] , \cur_error[11] , \cur_error[10] , 
        \cur_error[9] , \cur_error[8] , \cur_error[7] , \cur_error[6] , 
        \cur_error[5] , \cur_error[4] , \cur_error[3] , \cur_error[2] , 
        \cur_error[1] , \cur_error[0] }), .sr_prev({\sr_prev[12] , 
        \sr_prev[11] , \sr_prev[10] , \sr_prev[9] , \sr_prev[8] , 
        \sr_prev[7] , \sr_prev[6] , \sr_prev[5] , \sr_prev[4] , 
        \sr_prev[3] , \sr_prev[2] , \sr_prev[1] , \sr_prev[0] }), 
        .sr_new_0_0(\sr_new_0[12] ), .sr_new_1_0(\sr_new_1[12] ), 
        .int_enable(int_enable), .n_rst_c(n_rst_c), .clk_c(clk_c));
    controller_Z1_4 CONTROLLER (.state_0_d0(\state[1] ), .state_0_0(
        \state[0] ), .pwm_chg(pwm_chg), .sig_prev_0(sig_prev), 
        .sig_old_i_0_0(sig_old_i_0), .N_46_1(N_46_1), .avg_done(
        avg_done), .sig_old_i_0(sig_old_i_0_0), .sig_prev(sig_prev_0), 
        .sum_rdy(sum_rdy), .deriv_enable(deriv_enable), .calc_avg(
        calc_avg), .calc_int(calc_int), .pwm_enable(pwm_enable), 
        .sum_enable(sum_enable), .calc_error(calc_error), .avg_enable(
        avg_enable), .int_enable(int_enable), .pwm_chg_0(pwm_chg_0), 
        .avg_enable_0(avg_enable_0), .n_rst_c(n_rst_c), .clk_c(clk_c), 
        .avg_enable_1(avg_enable_1));
    sig_gen_0 FM_CYCLE (.primary_12_c(primary_12_c), .n_rst_c(n_rst_c), 
        .clk_c(clk_c), .sig_old_i_0(sig_old_i_0), .sig_prev(sig_prev));
    pid_sum_13s_4 SUM (.integral_i({\integral_i[25] , \integral_i[24] })
        , .integral({\integral[25] , \integral[24] , \integral[23] , 
        \integral[22] , \integral[21] , \integral[20] , \integral[19] , 
        \integral[18] , \integral[17] , \integral[16] , \integral[15] , 
        \integral[14] , \integral[13] , \integral[12] , \integral[11] , 
        \integral[10] , \integral[9] , \integral[8] , \integral[7] , 
        \integral[6] }), .sr_new({\sr_new[12] , \sr_new[11] , 
        \sr_new[10] , \sr_new[9] , \sr_new[8] , \sr_new[7] , 
        \sr_new[6] , \sr_new[5] , \sr_new[4] , \sr_new[3] , 
        \sr_new[2] , \sr_new[1] , \sr_new[0] }), .sr_new_0_0(
        \sr_new_0[12] ), .derivative_0(\derivative[12] ), .sr_new_1_0(
        \sr_new_1[12] ), .integral_0_0(\integral_0[25] ), 
        .integral_1_0(\integral_1[25] ), .sum_39(\sum[39] ), .sum_14(
        \sum[14] ), .sum_19(\sum[19] ), .sum_20(\sum[20] ), .sum_22(
        \sum[22] ), .sum_13(\sum[13] ), .sum_18(\sum[18] ), .sum_17(
        \sum[17] ), .sum_23(\sum[23] ), .sum_21(\sum[21] ), .sum_16(
        \sum[16] ), .sum_15(\sum[15] ), .sum_12(\sum[12] ), .sum_11(
        \sum[11] ), .sum_6(\sum[6] ), .sum_10(\sum[10] ), .sum_9(
        \sum[9] ), .sum_5(\sum[5] ), .sum_8(\sum[8] ), .sum_7(\sum[7] )
        , .sum_4(\sum[4] ), .sum_2_d0(\sum[2] ), .sum_1_d0(\sum[1] ), 
        .sum_0_d0(\sum[0] ), .sum_3(\sum[3] ), .sum_0_0(\sum_0[39] ), 
        .sum_1_0(\sum_1[39] ), .sum_2_0(\sum_2[39] ), .sum_enable(
        sum_enable), .sum_rdy(sum_rdy), .n_rst_c(n_rst_c), .clk_c(
        clk_c));
    sig_gen VD_SIG (.vd_done(vd_done), .n_rst_c(n_rst_c), .clk_c(clk_c)
        , .sig_old_i_0(sig_old_i_0_0), .sig_prev(sig_prev_0));
    spi_rx_12s_0 SPI (.cur_vd({\cur_vd[11] , \cur_vd[10] , \cur_vd[9] , 
        \cur_vd[8] , \cur_vd[7] , \cur_vd[6] , \cur_vd[5] , 
        \cur_vd[4] , \cur_vd[3] , \cur_vd[2] , \cur_vd[1] , 
        \cur_vd[0] }), .vd_done(vd_done), .cs_i_1_i(cs_i_1_i), 
        .cur_clk(cur_clk), .n_rst_c(n_rst_c), .din_12_c(din_12_c));
    integral_calc_13s_0_4 INTCALC (.sr_new({\sr_new[12] , \sr_new[11] , 
        \sr_new[10] , \sr_new[9] , \sr_new[8] , \sr_new[7] , 
        \sr_new[6] , \sr_new[5] , \sr_new[4] , \sr_new[3] , 
        \sr_new[2] , \sr_new[1] , \sr_new[0] }), .sr_old({\sr_old[12] , 
        \sr_old[11] , \sr_old[10] , \sr_old[9] , \sr_old[8] , 
        \sr_old[7] , \sr_old[6] , \sr_old[5] , \sr_old[4] , 
        \sr_old[3] , \sr_old[2] , \sr_old[1] , \sr_old[0] }), 
        .sr_new_1_0(\sr_new_1[12] ), .sr_new_0_0(\sr_new_0[12] ), 
        .integral({\integral[25] , \integral[24] , \integral[23] , 
        \integral[22] , \integral[21] , \integral[20] , \integral[19] , 
        \integral[18] , \integral[17] , \integral[16] , \integral[15] , 
        \integral[14] , \integral[13] , \integral[12] , \integral[11] , 
        \integral[10] , \integral[9] , \integral[8] , \integral[7] , 
        \integral[6] }), .integral_i({\integral_i[25] , 
        \integral_i[24] }), .integral_0_0(\integral_0[25] ), 
        .integral_1_0(\integral_1[25] ), .calc_int(calc_int), .N_46_1(
        N_46_1), .n_rst_c(n_rst_c), .clk_c(clk_c));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    error_calc_13s_12s_4 EC (.cur_error({\cur_error[12] , 
        \cur_error[11] , \cur_error[10] , \cur_error[9] , 
        \cur_error[8] , \cur_error[7] , \cur_error[6] , \cur_error[5] , 
        \cur_error[4] , \cur_error[3] , \cur_error[2] , \cur_error[1] , 
        \cur_error[0] }), .LED_12_i_0(\LED_12_i[5] ), .LED_12({
        \LED_12[7] , \LED_12[6] , LED_12[5], LED_12[4], LED_12[3], 
        LED_12[2], LED_12[1], LED_12[0]}), .average({\average[6] , 
        \average[5] , \average[4] , \average[3] , \average[2] }), 
        .calc_error(calc_error), .n_rst_c(n_rst_c), .clk_c(clk_c));
    derivative_calc_13s_4 DCALC (.derivative_0(\derivative[12] ), 
        .sr_prev({\sr_prev[12] , \sr_prev[11] , \sr_prev[10] , 
        \sr_prev[9] , \sr_prev[8] , \sr_prev[7] , \sr_prev[6] , 
        \sr_prev[5] , \sr_prev[4] , \sr_prev[3] , \sr_prev[2] , 
        \sr_prev[1] , \sr_prev[0] }), .sr_new({\sr_new[11] , 
        \sr_new[10] , \sr_new[9] , \sr_new[8] , \sr_new[7] , 
        \sr_new[6] , \sr_new[5] , \sr_new[4] , \sr_new[3] , 
        \sr_new[2] , \sr_new[1] , \sr_new[0] }), .sr_new_0_0(
        \sr_new_0[12] ), .deriv_enable(deriv_enable), .n_rst_c(n_rst_c)
        , .clk_c(clk_c));
    pwm_tx_200s_32s_13s_10_216s_51s PWM_TX (.off_div({\off_div[31] , 
        \off_div[30] , \off_div[29] , \off_div[28] , \off_div[27] , 
        \off_div[26] , \off_div[25] , \off_div[24] , \off_div[23] , 
        \off_div[22] , \off_div[21] , \off_div[20] , \off_div[19] , 
        \off_div[18] , \off_div[17] , \off_div[16] , \off_div[15] , 
        \off_div[14] , \off_div[13] , \off_div[12] , \off_div[11] , 
        \off_div[10] , \off_div[9] , \off_div[8] , \off_div[7] , 
        \off_div[6] , \off_div[5] , \off_div[4] , \off_div[3] , 
        \off_div[2] , \off_div[1] , \off_div[0] }), .act_ctl_5_i(
        act_ctl_5_i), .act_ctl_5_0(act_ctl_5_0), .act_ctl_5_8(
        act_ctl_5_8), .pwm_chg(pwm_chg), .pwm_chg_0(pwm_chg_0), 
        .n_rst_c(n_rst_c), .clk_c(clk_c), .act_ctl_5(act_ctl_5), 
        .act_ctl_5_9(act_ctl_5_9), .act_ctl_5_4(act_ctl_5_4), 
        .act_ctl_5_3(act_ctl_5_3), .act_ctl_5_7(act_ctl_5_7), 
        .primary_12_c(primary_12_c));
    spi_clk_11s_0 SPICLK (.cur_clk(cur_clk), .n_rst_c(n_rst_c), .clk_c(
        clk_c));
    
endmodule


module pwm_ctl_200s_32s_13s_0_1_2_2(
       sum_8,
       sum_39,
       sum_10,
       sum_11,
       sum_12,
       sum_13,
       sum_15,
       sum_16,
       sum_17,
       sum_18,
       sum_19,
       sum_20,
       sum_21,
       sum_22,
       sum_23,
       sum_14,
       sum_9,
       sum_2_d0,
       sum_1_d0,
       sum_0_d0,
       sum_7,
       sum_6,
       sum_4,
       sum_3,
       sum_5,
       off_div,
       sum_1_0,
       sum_0_0,
       sum_2_0,
       n_rst_c,
       clk_c,
       pwm_enable,
       pwm_rdy
    );
input  sum_8;
input  sum_39;
input  sum_10;
input  sum_11;
input  sum_12;
input  sum_13;
input  sum_15;
input  sum_16;
input  sum_17;
input  sum_18;
input  sum_19;
input  sum_20;
input  sum_21;
input  sum_22;
input  sum_23;
input  sum_14;
input  sum_9;
input  sum_2_d0;
input  sum_1_d0;
input  sum_0_d0;
input  sum_7;
input  sum_6;
input  sum_4;
input  sum_3;
input  sum_5;
output [31:0] off_div;
input  sum_1_0;
input  sum_0_0;
input  sum_2_0;
input  n_rst_c;
input  clk_c;
input  pwm_enable;
output pwm_rdy;

    wire un1_state_2_0, un5lt31, next_off_div_2_sqmuxa_11, 
        \state[1]_net_1 , \state_d_0[2] , \state[0]_net_1 , N_16, 
        \DWACT_FINC_E[4] , N_13, \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , 
        ADD_32x32_fast_I321_Y_0, ADD_32x32_fast_I258_Y_3, N625, N610, 
        ADD_32x32_fast_I258_Y_2, N551, N544, ADD_32x32_fast_I258_Y_1, 
        N479, N482, ADD_32x32_fast_I258_Y_0, ADD_32x32_fast_I320_Y_0, 
        ADD_32x32_fast_I313_Y_0, ADD_32x32_fast_I259_Y_3, N627, N612, 
        ADD_32x32_fast_I259_Y_2, N553, N546, ADD_32x32_fast_I259_Y_1, 
        N481, N484, ADD_32x32_fast_I259_Y_0, 
        ADD_32x32_fast_I258_un1_Y_0, N626, ADD_32x32_fast_I318_Y_0, 
        ADD_32x32_fast_I319_Y_0, ADD_32x32_fast_I317_Y_0, 
        ADD_32x32_fast_I314_Y_0, ADD_32x32_fast_I315_Y_0, 
        ADD_32x32_fast_I316_Y_0, ADD_32x32_fast_I266_Y_0, N641, 
        ADD_32x32_fast_I260_Y_2, N614, N629, ADD_32x32_fast_I260_Y_1, 
        I158_un1_Y, I98_un1_Y, ADD_32x32_fast_I261_Y_2, N616, N631, 
        ADD_32x32_fast_I261_Y_1, N557, N550, ADD_32x32_fast_I261_Y_0, 
        I100_un1_Y, ADD_32x32_fast_I312_Y_0, ADD_32x32_fast_I304_Y_0, 
        \un1_sum_adj[14] , ADD_32x32_fast_I259_un1_Y_0, N628, 
        ADD_32x32_fast_I262_Y_1, N618, N633, ADD_32x32_fast_I262_Y_0, 
        I162_un1_Y, ADD_32x32_fast_I310_Y_0, ADD_32x32_fast_I311_Y_0, 
        ADD_32x32_fast_I309_Y_0, ADD_32x32_fast_I266_un1_Y_0, N642, 
        ADD_32x32_fast_I265_Y_1, N639, N624, ADD_32x32_fast_I265_Y_0, 
        N565, N558, ADD_32x32_fast_I263_Y_1, N635, N620, 
        ADD_32x32_fast_I263_Y_0, N561, N554, ADD_32x32_fast_I264_Y_1, 
        N622, N637, ADD_32x32_fast_I264_Y_0, N556, N563, N555, 
        ADD_32x32_fast_I306_Y_0, ADD_32x32_fast_I308_Y_0, 
        ADD_32x32_fast_I307_Y_0, ADD_32x32_fast_I302_Y_0, 
        \un1_sum_adj[12] , ADD_32x32_fast_I303_Y_0, 
        \sum_adj[21]_net_1 , ADD_32x32_fast_I260_un1_Y_0, N630, 
        ADD_32x32_fast_I261_un1_Y_0, N632, ADD_32x32_fast_I301_Y_0, 
        \sum_adj[19]_net_1 , ADD_32x32_fast_I262_un1_Y_0, N634, 
        ADD_32x32_fast_I269_Y_0, N647, ADD_32x32_fast_I270_Y_0, N649, 
        ADD_32x32_fast_I298_Y_0, \un1_sum_adj[8] , 
        ADD_32x32_fast_I299_Y_0, \un1_sum_adj[9] , 
        ADD_32x32_fast_I300_Y_0, \sum_adj_RNIJIDD[18]_net_1 , 
        ADD_32x32_fast_I263_un1_Y_0, N636, ADD_32x32_fast_I265_un1_Y_0, 
        N640, ADD_32x32_fast_I264_un1_Y_0, N638, 
        ADD_32x32_fast_I296_Y_0, \sum_adj[14]_net_1 , 
        ADD_32x32_fast_I271_Y_0, ADD_32x32_fast_I271_un1_Y_0, 
        ADD_32x32_fast_I272_Y_0, ADD_32x32_fast_I272_un1_Y_0, 
        ADD_32x32_fast_I295_Y_0, \un1_sum_adj[5] , 
        ADD_32x32_fast_I294_Y_0, \un1_sum_adj[4] , 
        ADD_32x32_fast_I268_un1_Y_0, N646, ADD_32x32_fast_I293_Y_0, 
        \sum_adj[11]_net_1 , N586, N594, N601, N538, N654, 
        ADD_32x32_fast_I292_Y_0, \sum_adj[10]_net_1 , 
        next_off_div_2_sqmuxa_9, next_off_div_2_sqmuxa_8, 
        next_off_div16, un1_off_divlto31_9, next_off_div_2_sqmuxa_0, 
        next_off_div_2_sqmuxa_7, next_off_div_2_sqmuxa_5, 
        next_off_div_2_sqmuxa_3, ADD_32x32_fast_I291_Y_0, 
        \un1_sum_adj[1] , un5lto20_2, un5lto20_1, un5lto14_2, 
        un5lto14_1, un1_off_divlto31_22, un1_off_divlto31_15, 
        un1_off_divlto31_14, un1_off_divlto31_20, un1_off_divlto31_21, 
        un1_off_divlto31_13, un1_off_divlto31_12, un1_off_divlto31_17, 
        un1_off_divlto31_10, un1_off_divlt31, un1_off_divlto31_0, 
        un5lto9, un1_off_divlto31_8, un1_off_divlto31_6, 
        un1_off_divlto31_4, un1_off_divlto31_2, un5lto7_1, N483, N487, 
        un5lt9, un5lto4, un5lt4, N751, N784, I262_un1_Y, N793, 
        I267_un1_Y, N644, N659, \un1_off_div_1[27] , 
        \un1_off_div_1[15] , \un1_sum_adj[15] , N781, N767, I228_un1_Y, 
        \un1_off_div_1[5] , N661, N779, I273_un1_Y, I240_un1_Y, N656, 
        \sum_adj_RNIH9EC[8]_net_1 , N749, N761, N799, 
        \un1_off_div_1[0] , next_off_div_1_sqmuxa, N753, N787, 
        I270_un1_Y, N650, N599, \un1_off_div_1[19] , N759, N796, N769, 
        I230_un1_Y, I268_un1_Y, \un1_off_div_1[20] , I269_un1_Y, N648, 
        N663, N765, N657, un5lt16, \un1_off_div_1[3] , N755, N790, 
        N763, N802, \un1_off_div_1[10] , \un1_off_div_1[17] , 
        I238_un1_Y, \un1_off_div_1[18] , I236_un1_Y, 
        \un1_off_div_1[7] , \un1_sum_adj[7] , \next_off_div[4] , N395, 
        N396, N485, N651, N653, \nsum_adj_5[8] , I_23_11, 
        \nsum_adj_5[10] , I_28_3, \nsum_adj_5[11] , I_32_3, 
        \nsum_adj_5[12] , I_35_3, \nsum_adj_5[13] , I_37_3, 
        \nsum_adj_5[15] , I_43_3, \nsum_adj_5[16] , I_46_3, 
        \nsum_adj_5[17] , I_49_3, \nsum_adj_5[18] , I_53_3, 
        \nsum_adj_5[19] , I_56_3, \nsum_adj_5[20] , I_59_3, 
        \nsum_adj_5[21] , I_62_3, \nsum_adj_5[22] , I_65_3, 
        \nsum_adj_5[23] , I_70_3, \sum_adj[12]_net_1 , 
        \next_off_div[18] , \state_d[2] , \next_off_div[17] , 
        \next_off_div[7] , state_176_d, \next_off_div[10] , 
        \next_off_div[24] , \next_off_div[28] , 
        \state_RNI51T1I_0[1]_net_1 , \next_off_div[3] , un5lt14, 
        \next_off_div[11] , \next_off_div[23] , \next_off_div[20] , 
        \next_off_div[21] , N645, \next_off_div[26] , 
        \next_off_div[19] , N486, N564, N571, \next_off_div[29] , 
        \next_off_div[0] , \next_off_div[25] , I247_un1_Y, 
        \nsum_adj_5[14] , I_40_3, \nsum_adj_5[9] , I_26_3, 
        \next_off_div[2] , \next_off_div[1] , \next_off_div[16] , 
        \next_off_div[31] , N552, N573, N566, N655, \next_off_div[5] , 
        \next_off_div[22] , N562, \next_off_div[15] , 
        \sum_adj[23]_net_1 , I246_un1_Y, N643, N429, N428, 
        \next_off_div[30] , \next_off_div[27] , \state_ns[0] , N_311_i, 
        \next_off_div[8] , \next_off_div[9] , \next_off_div[12] , 
        \next_off_div[13] , \next_off_div[14] , N383, N392, N393, N401, 
        N402, N404, N408, N521, N522, N407, N523, N524, N525, N532, 
        N389, N533, N390, N534, N386, N537, N387, \sum_adj[8]_net_1 , 
        N580, N519, N515, N584, N587, N526, N589, N528, N590, N529, 
        N591, N530, N527, N593, N597, N536, N598, I150_un1_Y, N535, 
        N572, N576, N592, N579, N518, N514, N417, N511, N507, N510, 
        N506, N414, N410, N413, N416, N419, N422, N423, N425, N426, 
        N513, N516, N517, N520, N489, N575, N578, N581, N582, N583, 
        N585, N569, N568, N567, N570, \sum_adj[22]_net_1 , 
        \sum_adj[20]_net_1 , \sum_adj[18]_net_1 , \sum_adj[17]_net_1 , 
        \sum_adj[16]_net_1 , \sum_adj[15]_net_1 , I196_un1_Y, 
        I204_un1_Y, N595, N596, N588, I190_un1_Y, N531, N398, N503, 
        N502, \next_off_div[6] , N490, N498, N499, N497, N493, N560, 
        N495, N491, N492, N494, N496, \sum_adj[9]_net_1 , N500, N501, 
        N504, N505, N432, N508, N509, \sum_adj[13]_net_1 , N577, N574, 
        N512, N_2, \DWACT_FINC_E[29] , \DWACT_FINC_E[13] , 
        \DWACT_FINC_E[33] , \DWACT_FINC_E[34] , \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[5] , \DWACT_FINC_E[15] , N_3, \DWACT_FINC_E[28] , 
        \DWACT_FINC_E[16] , N_4, N_5, \DWACT_FINC_E[14] , N_6, 
        \DWACT_FINC_E[9] , \DWACT_FINC_E[12] , N_7, \DWACT_FINC_E[10] , 
        \DWACT_FINC_E[0] , N_8, \DWACT_FINC_E[11] , N_9, N_10, N_11, 
        \DWACT_FINC_E[8] , N_12, N_14, N_15, \DWACT_FINC_E[3] , N_17, 
        GND, VCC;
    
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I59_Y (.A(sum_2_0), .B(
        off_div[17]), .C(N432), .Y(N505));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_2 (.A(N551), .B(N544), 
        .C(ADD_32x32_fast_I258_Y_1), .Y(ADD_32x32_fast_I258_Y_2));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I10_P0N (.A(
        \sum_adj_RNIJIDD[18]_net_1 ), .B(off_div[10]), .Y(N414));
    DFN1C0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[0]_net_1 ));
    DFN1E0C0 \off_div[29]  (.D(\next_off_div[29] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[29]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y_0 (.A(N556), .B(N563), 
        .C(N555), .Y(ADD_32x32_fast_I264_Y_0));
    DFN1E0C0 \off_div[26]  (.D(\next_off_div[26] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[26]));
    XNOR2 un1_nsum_adj_I_43 (.A(sum_15), .B(N_10), .Y(I_43_3));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I247_Y (.A(I247_un1_Y), .B(
        N651), .Y(N796));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I108_Y (.A(N496), .B(N492), 
        .Y(N557));
    AND3 un1_nsum_adj_I_48 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[11] ), .Y(N_8));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I47_Y (.A(off_div[23]), .B(
        off_div[22]), .C(sum_1_0), .Y(N493));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I3_P0N (.A(sum_1_0), .B(
        \sum_adj[11]_net_1 ), .C(off_div[3]), .Y(N393));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I165_Y (.A(N562), .B(N554), 
        .Y(N620));
    DFN1E0C0 \off_div[31]  (.D(\next_off_div[31] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[31]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I149_Y (.A(N537), .B(N533), 
        .Y(N598));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I135_Y (.A(N523), .B(N519), 
        .Y(N584));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I147_Y (.A(N535), .B(N531), 
        .Y(N596));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I121_Y (.A(N505), .B(N509), 
        .Y(N570));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I272_Y_0 (.A(
        ADD_32x32_fast_I272_un1_Y_0), .B(N638), .C(N637), .Y(
        ADD_32x32_fast_I272_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I173_Y (.A(N562), .B(N570), 
        .Y(N628));
    MX2 \sum_adj_RNO[9]  (.A(sum_9), .B(I_26_3), .S(sum_0_0), .Y(
        \nsum_adj_5[9] ));
    XA1 \off_div_RNO[22]  (.A(N767), .B(ADD_32x32_fast_I312_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[22] ));
    NOR2A \off_div_RNIH86K[29]  (.A(\state[0]_net_1 ), .B(off_div[29]), 
        .Y(next_off_div_2_sqmuxa_5));
    DFN1E1C0 \sum_adj[23]  (.D(\nsum_adj_5[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[23]_net_1 ));
    OA1 \off_div_RNI4R23[1]  (.A(un5lto4), .B(un5lt4), .C(un5lto7_1), 
        .Y(un5lt9));
    NOR3 un1_nsum_adj_I_41 (.A(sum_13), .B(sum_12), .C(sum_14), .Y(
        \DWACT_FINC_E[9] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I203_Y (.A(N594), .B(N601), 
        .C(N593), .Y(N659));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I155_Y (.A(N552), .B(N544), 
        .Y(N610));
    NOR2B un1_nsum_adj_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_13));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I86_Y (.A(N389), .B(N393), .C(
        N392), .Y(N532));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I200_Y (.A(N597), .B(N590), 
        .C(N589), .Y(N655));
    XNOR2 un1_nsum_adj_I_37 (.A(sum_13), .B(N_12), .Y(I_37_3));
    MX2 \sum_adj_RNO[15]  (.A(sum_15), .B(I_43_3), .S(sum_0_0), .Y(
        \nsum_adj_5[15] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I315_Y_0 (.A(off_div[25]), 
        .B(sum_39), .Y(ADD_32x32_fast_I315_Y_0));
    NOR3 un1_nsum_adj_I_10 (.A(sum_2_d0), .B(sum_1_d0), .C(sum_0_d0), 
        .Y(\DWACT_FINC_E[0] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I84_Y (.A(N392), .B(N396), .C(
        N395), .Y(N530));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I130_Y (.A(N518), .B(N515), 
        .C(N514), .Y(N579));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I266_Y (.A(
        ADD_32x32_fast_I266_un1_Y_0), .B(N657), .C(
        ADD_32x32_fast_I266_Y_0), .Y(N765));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I118_Y (.A(N506), .B(N503), 
        .C(N502), .Y(N567));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I69_Y (.A(off_div[12]), .B(
        \un1_sum_adj[12] ), .C(N417), .Y(N515));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I262_Y_0 (.A(N551), .B(
        I162_un1_Y), .Y(ADD_32x32_fast_I262_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I202_Y (.A(N592), .B(N599), 
        .C(N591), .Y(N657));
    MX2 \sum_adj_RNO[16]  (.A(sum_16), .B(I_46_3), .S(sum_0_0), .Y(
        \nsum_adj_5[16] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I309_Y_0 (.A(off_div[19]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I309_Y_0));
    NOR3A \off_div_RNIG5HD1[30]  (.A(next_off_div_2_sqmuxa_5), .B(
        off_div[30]), .C(off_div[28]), .Y(next_off_div_2_sqmuxa_8));
    MX2 \off_div_RNO[3]  (.A(next_off_div16), .B(\un1_off_div_1[3] ), 
        .S(\state_d_0[2] ), .Y(\next_off_div[3] ));
    XNOR2 un1_nsum_adj_I_70 (.A(sum_23), .B(N_2), .Y(I_70_3));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I76_Y (.A(N404), .B(N408), .C(
        N407), .Y(N522));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I4_G0N (.A(\un1_sum_adj[4] )
        , .B(off_div[4]), .Y(N395));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I1_P0N (.A(\un1_sum_adj[1] ), 
        .B(off_div[1]), .Y(N387));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I13_G0N (.A(sum_0_0), .B(
        \sum_adj[21]_net_1 ), .C(off_div[13]), .Y(N422));
    DFN1E0C0 \off_div[15]  (.D(\next_off_div[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[15]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I150_Y (.A(I150_un1_Y), .B(
        N534), .Y(N599));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I144_Y (.A(N532), .B(N529), 
        .C(N528), .Y(N593));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I74_Y (.A(N407), .B(
        off_div[9]), .C(\un1_sum_adj[9] ), .Y(N520));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I50_Y (.A(off_div[21]), .B(
        off_div[20]), .C(sum_2_0), .Y(N496));
    DFN1E0C0 \off_div[13]  (.D(\next_off_div[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[13]));
    XNOR2 un1_nsum_adj_I_62 (.A(sum_21), .B(N_4), .Y(I_62_3));
    MX2 \sum_adj_RNO[20]  (.A(sum_20), .B(I_59_3), .S(sum_0_0), .Y(
        \nsum_adj_5[20] ));
    NOR3C \off_div_RNI1OGI1[17]  (.A(off_div[18]), .B(off_div[17]), .C(
        un5lto20_1), .Y(un5lto20_2));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I293_Y_0 (.A(sum_0_0), .B(
        \sum_adj[11]_net_1 ), .C(off_div[3]), .Y(
        ADD_32x32_fast_I293_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I272_un1_Y_0 (.A(N538), .B(
        N654), .Y(ADD_32x32_fast_I272_un1_Y_0));
    NOR2B \off_div_RNIUP8P[19]  (.A(off_div[20]), .B(off_div[19]), .Y(
        un5lto20_1));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I319_Y_0 (.A(off_div[29]), 
        .B(sum_39), .Y(ADD_32x32_fast_I319_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I265_Y_0 (.A(N565), .B(N558), 
        .C(N557), .Y(ADD_32x32_fast_I265_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I179_Y (.A(N568), .B(N576), 
        .Y(N634));
    XA1 \off_div_RNO[24]  (.A(N763), .B(ADD_32x32_fast_I314_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[24] ));
    XNOR2 un1_nsum_adj_I_35 (.A(sum_12), .B(N_13), .Y(I_35_3));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I309_Y (.A(I270_un1_Y), .B(
        ADD_32x32_fast_I270_Y_0), .C(ADD_32x32_fast_I309_Y_0), .Y(
        \un1_off_div_1[19] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I177_Y (.A(N566), .B(N574), 
        .Y(N632));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I51_Y (.A(off_div[20]), .B(
        off_div[21]), .C(sum_2_0), .Y(N497));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I308_Y_0 (.A(off_div[18]), 
        .B(sum_39), .Y(ADD_32x32_fast_I308_Y_0));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I2_P0N (.A(sum_0_0), .B(
        \sum_adj[10]_net_1 ), .C(off_div[2]), .Y(N390));
    DFN1E0P0 \off_div[7]  (.D(\next_off_div[7] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[7]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I196_Y (.A(I196_un1_Y), .B(
        N585), .Y(N651));
    AO1C \state_RNI51T1I_0[1]  (.A(un5lt31), .B(
        next_off_div_2_sqmuxa_11), .C(\state[1]_net_1 ), .Y(
        \state_RNI51T1I_0[1]_net_1 ));
    AND3 un1_nsum_adj_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[6] ));
    XOR2 \sum_adj_RNIROSJ[20]  (.A(\sum_adj[20]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[12] ));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I268_Y (.A(I230_un1_Y), .B(
        N629), .C(I268_un1_Y), .Y(N769));
    OA1 \off_div_RNIHJFG[10]  (.A(un5lto9), .B(un5lt9), .C(off_div[10])
        , .Y(un5lt14));
    DFN1E0C0 \off_div[9]  (.D(\next_off_div[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[9]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I37_Y (.A(off_div[27]), .B(
        off_div[28]), .C(sum_1_0), .Y(N483));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_1 (.A(N481), .B(N484), 
        .C(ADD_32x32_fast_I259_Y_0), .Y(ADD_32x32_fast_I259_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I186_Y (.A(N583), .B(N576), 
        .C(N575), .Y(N641));
    DFN1E0C0 \off_div[11]  (.D(\next_off_div[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[11]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I145_Y (.A(N529), .B(N533), 
        .Y(N594));
    NOR2A un1_nsum_adj_I_63 (.A(\DWACT_FINC_E[15] ), .B(sum_21), .Y(
        \DWACT_FINC_E[16] ));
    DFN1E1C0 \sum_adj[18]  (.D(\nsum_adj_5[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[18]_net_1 ));
    MX2 un1_off_div_1_0_0_ADD_32x32_fast_I92_Y (.A(sum_0_0), .B(
        off_div[0]), .S(\sum_adj[8]_net_1 ), .Y(N538));
    AND3 un1_nsum_adj_I_68 (.A(\DWACT_FINC_E[34] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[29] ));
    XA1 \off_div_RNO[13]  (.A(N787), .B(ADD_32x32_fast_I303_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[13] ));
    MX2 \sum_adj_RNO[21]  (.A(sum_21), .B(I_62_3), .S(sum_0_0), .Y(
        \nsum_adj_5[21] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I318_Y_0 (.A(off_div[28]), 
        .B(sum_39), .Y(ADD_32x32_fast_I318_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I191_Y (.A(N588), .B(N580), 
        .Y(N646));
    MX2 \sum_adj_RNO[22]  (.A(sum_22), .B(I_65_3), .S(sum_1_0), .Y(
        \nsum_adj_5[22] ));
    MX2 \off_div_RNO[15]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[15] ), .S(\state_d[2] ), .Y(\next_off_div[15] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y (.A(
        ADD_32x32_fast_I258_un1_Y_0), .B(N781), .C(
        ADD_32x32_fast_I258_Y_3), .Y(N749));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I14_P0N (.A(\un1_sum_adj[14] )
        , .B(off_div[14]), .Y(N426));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I122_Y (.A(N510), .B(N507), 
        .C(N506), .Y(N571));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I89_Y (.A(N387), .B(N390), 
        .Y(N535));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I262_Y_1 (.A(N618), .B(N633), 
        .C(ADD_32x32_fast_I262_Y_0), .Y(ADD_32x32_fast_I262_Y_1));
    AND2 un1_nsum_adj_I_44 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[9] ), .Y(\DWACT_FINC_E[10] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I265_Y (.A(
        ADD_32x32_fast_I265_un1_Y_0), .B(N802), .C(
        ADD_32x32_fast_I265_Y_1), .Y(N763));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I181_Y (.A(N570), .B(N578), 
        .Y(N636));
    AND3 un1_nsum_adj_I_61 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[15] ), .Y(N_4));
    NOR2 un1_nsum_adj_I_47 (.A(sum_16), .B(sum_15), .Y(
        \DWACT_FINC_E[11] ));
    DFN1E1C0 \sum_adj[9]  (.D(\nsum_adj_5[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[9]_net_1 ));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I60_Y (.A(N428), .B(sum_2_0), 
        .C(off_div[16]), .Y(N506));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I4_P0N (.A(\un1_sum_adj[4] ), 
        .B(off_div[4]), .Y(N396));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I307_Y (.A(I238_un1_Y), .B(
        ADD_32x32_fast_I272_Y_0), .C(ADD_32x32_fast_I307_Y_0), .Y(
        \un1_off_div_1[17] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I174_Y (.A(N564), .B(N571), 
        .C(N563), .Y(N629));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I140_Y (.A(N528), .B(N525), 
        .C(N524), .Y(N589));
    DFN1E1C0 \sum_adj[11]  (.D(\nsum_adj_5[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[11]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y_1 (.A(N635), .B(N620), 
        .C(ADD_32x32_fast_I263_Y_0), .Y(ADD_32x32_fast_I263_Y_1));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I246_Y (.A(I246_un1_Y), .B(
        N649), .Y(N793));
    NOR2B \off_div_RNO[27]  (.A(\un1_off_div_1[27] ), .B(\state_d[2] ), 
        .Y(\next_off_div[27] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I291_Y_0 (.A(off_div[1]), .B(
        \un1_sum_adj[1] ), .Y(ADD_32x32_fast_I291_Y_0));
    NOR3B un1_nsum_adj_I_36 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .C(sum_12), .Y(N_12));
    NOR3C \off_div_RNIT951[6]  (.A(off_div[6]), .B(off_div[7]), .C(
        off_div[5]), .Y(un5lto7_1));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I13_P0N (.A(sum_0_0), .B(
        \sum_adj[21]_net_1 ), .C(off_div[13]), .Y(N423));
    DFN1E0C0 \off_div[25]  (.D(\next_off_div[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[25]));
    XA1 \off_div_RNO[1]  (.A(N538), .B(ADD_32x32_fast_I291_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[1] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I61_Y (.A(N429), .B(N432), 
        .Y(N507));
    DFN1E1C0 \sum_adj[22]  (.D(\nsum_adj_5[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[22]_net_1 ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I79_Y (.A(off_div[7]), .B(
        \un1_sum_adj[7] ), .C(N402), .Y(N525));
    NOR2 \off_div_RNIPMAP[31]  (.A(off_div[31]), .B(off_div[21]), .Y(
        next_off_div_2_sqmuxa_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I150_un1_Y (.A(N535), .B(
        N538), .Y(I150_un1_Y));
    OA1 \off_div_RNIEQ41[1]  (.A(off_div[0]), .B(off_div[1]), .C(
        off_div[2]), .Y(un5lt4));
    DFN1E0C0 \off_div[23]  (.D(\next_off_div[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[23]));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I304_Y_0 (.A(off_div[14]), 
        .B(\un1_sum_adj[14] ), .Y(ADD_32x32_fast_I304_Y_0));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I298_Y_0 (.A(off_div[8]), .B(
        \un1_sum_adj[8] ), .Y(ADD_32x32_fast_I298_Y_0));
    XA1 \off_div_RNO[9]  (.A(N799), .B(ADD_32x32_fast_I299_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[9] ));
    NOR2 \off_div_RNITN7P[14]  (.A(off_div[14]), .B(off_div[15]), .Y(
        un1_off_divlto31_6));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y_1 (.A(N622), .B(N637), 
        .C(ADD_32x32_fast_I264_Y_0), .Y(ADD_32x32_fast_I264_Y_1));
    GND GND_i (.Y(GND));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I95_Y (.A(N479), .B(N483), 
        .Y(N544));
    DFN1E1C0 \sum_adj[14]  (.D(\nsum_adj_5[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[14]_net_1 ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I98_un1_Y (.A(N486), .B(
        N483), .Y(I98_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I138_Y (.A(N526), .B(N523), 
        .C(N522), .Y(N587));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y (.A(
        ADD_32x32_fast_I259_un1_Y_0), .B(N784), .C(
        ADD_32x32_fast_I259_Y_3), .Y(N751));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I43_Y (.A(off_div[24]), .B(
        off_div[25]), .C(sum_1_0), .Y(N489));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I123_Y (.A(N507), .B(N511), 
        .Y(N572));
    NOR3B \state_RNIP9T79[1]  (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .C(next_off_div16), .Y(
        next_off_div_1_sqmuxa));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I175_Y (.A(N564), .B(N572), 
        .Y(N630));
    NOR3B un1_nsum_adj_I_45 (.A(\DWACT_FINC_E[10] ), .B(
        \DWACT_FINC_E[6] ), .C(sum_15), .Y(N_9));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I106_Y (.A(N490), .B(N494), 
        .Y(N555));
    MX2 \sum_adj_RNO[10]  (.A(sum_10), .B(I_28_3), .S(sum_0_0), .Y(
        \nsum_adj_5[10] ));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I317_Y (.A(I262_un1_Y), .B(
        ADD_32x32_fast_I262_Y_1), .C(ADD_32x32_fast_I317_Y_0), .Y(
        \un1_off_div_1[27] ));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I11_G0N (.A(sum_1_0), .B(
        \sum_adj[19]_net_1 ), .C(off_div[11]), .Y(N416));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I314_Y_0 (.A(off_div[24]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I314_Y_0));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I271_un1_Y_0 (.A(N586), .B(
        N594), .C(N601), .Y(ADD_32x32_fast_I271_un1_Y_0));
    DFN1E0C0 \off_div[21]  (.D(\next_off_div[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[21]));
    XA1B \off_div_RNO[11]  (.A(N793), .B(ADD_32x32_fast_I301_Y_0), .C(
        \state[0]_net_1 ), .Y(\next_off_div[11] ));
    XNOR2 un1_nsum_adj_I_40 (.A(sum_14), .B(N_11), .Y(I_40_3));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I42_Y (.A(off_div[25]), .B(
        off_div[24]), .C(sum_1_0), .Y(I100_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y (.A(
        ADD_32x32_fast_I263_un1_Y_0), .B(N796), .C(
        ADD_32x32_fast_I263_Y_1), .Y(N759));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I248_Y (.A(N654), .B(N538), 
        .C(N653), .Y(N799));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I301_Y_0 (.A(sum_2_0), .B(
        \sum_adj[19]_net_1 ), .C(off_div[11]), .Y(
        ADD_32x32_fast_I301_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y (.A(
        ADD_32x32_fast_I260_un1_Y_0), .B(N787), .C(
        ADD_32x32_fast_I260_Y_2), .Y(N753));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I306_Y_0 (.A(off_div[16]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I306_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I80_Y (.A(N398), .B(N402), .C(
        N401), .Y(N526));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I101_Y (.A(N489), .B(N485), 
        .Y(N550));
    DFN1E1C0 \sum_adj[13]  (.D(\nsum_adj_5[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[13]_net_1 ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I265_un1_Y_0 (.A(N624), .B(
        N640), .Y(ADD_32x32_fast_I265_un1_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I170_Y (.A(N567), .B(N560), 
        .C(I162_un1_Y), .Y(N625));
    DFN1E0C0 \off_div[5]  (.D(\next_off_div[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[5]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I7_G0N (.A(\un1_sum_adj[7] )
        , .B(off_div[7]), .Y(N404));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I57_Y (.A(off_div[18]), .B(
        off_div[17]), .C(sum_2_0), .Y(N503));
    XOR2 \state_RNO[1]  (.A(\state[1]_net_1 ), .B(\state[0]_net_1 ), 
        .Y(N_311_i));
    NOR2A \state_RNIRC2F_0[1]  (.A(\state[1]_net_1 ), .B(
        \state[0]_net_1 ), .Y(\state_d[2] ));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I308_Y (.A(I236_un1_Y), .B(
        ADD_32x32_fast_I271_Y_0), .C(ADD_32x32_fast_I308_Y_0), .Y(
        \un1_off_div_1[18] ));
    MX2 \sum_adj_RNO[11]  (.A(sum_11), .B(I_32_3), .S(sum_0_0), .Y(
        \nsum_adj_5[11] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I321_Y_0 (.A(off_div[31]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I321_Y_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I116_Y (.A(N500), .B(N504), 
        .Y(N565));
    NOR3C \off_div_RNIPFSO4[16]  (.A(un1_off_divlto31_15), .B(
        un1_off_divlto31_14), .C(un1_off_divlto31_20), .Y(
        un1_off_divlto31_22));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I311_Y_0 (.A(off_div[21]), 
        .B(sum_39), .Y(ADD_32x32_fast_I311_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I269_Y_0 (.A(N647), .B(N632), 
        .C(N631), .Y(ADD_32x32_fast_I269_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I81_Y (.A(off_div[5]), .B(
        \un1_sum_adj[5] ), .C(N402), .Y(N527));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I245_Y (.A(N648), .B(N663), 
        .C(N647), .Y(N790));
    MX2 \sum_adj_RNO[12]  (.A(sum_12), .B(I_35_3), .S(sum_0_0), .Y(
        \nsum_adj_5[12] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I316_Y_0 (.A(off_div[26]), 
        .B(sum_39), .Y(ADD_32x32_fast_I316_Y_0));
    AND3 un1_nsum_adj_I_64 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[16] ), .Y(N_3));
    NOR3 un1_nsum_adj_I_67 (.A(sum_2_d0), .B(sum_1_d0), .C(sum_0_d0), 
        .Y(\DWACT_FINC_E[34] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I70_Y (.A(N413), .B(N417), .C(
        N416), .Y(N516));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I192_Y (.A(N589), .B(N582), 
        .C(N581), .Y(N647));
    DFN1E0C0 \off_div[30]  (.D(\next_off_div[30] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[30]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I265_Y_1 (.A(N639), .B(N624), 
        .C(ADD_32x32_fast_I265_Y_0), .Y(ADD_32x32_fast_I265_Y_1));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I129_Y (.A(N513), .B(N517), 
        .Y(N578));
    XNOR2 un1_nsum_adj_I_46 (.A(sum_16), .B(N_9), .Y(I_46_3));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I182_Y (.A(N579), .B(N572), 
        .C(N571), .Y(N637));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I127_Y (.A(N511), .B(N515), 
        .Y(N576));
    AND3 un1_nsum_adj_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_17));
    VCC VCC_i (.Y(VCC));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I249_Y (.A(N656), .B(
        \sum_adj_RNIH9EC[8]_net_1 ), .C(N655), .Y(N802));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I0_G0N (.A(off_div[0]), .B(
        sum_39), .Y(N383));
    AND3 un1_nsum_adj_I_39 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[8] ), .Y(N_11));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I196_un1_Y (.A(N593), .B(
        N586), .Y(I196_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I45_Y (.A(off_div[24]), .B(
        off_div[23]), .C(sum_1_0), .Y(N491));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I111_Y (.A(N499), .B(N495), 
        .Y(N560));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I71_Y (.A(N414), .B(N417), 
        .Y(N517));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I9_G0N (.A(\un1_sum_adj[9] )
        , .B(off_div[9]), .Y(N410));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I228_un1_Y (.A(N643), .B(
        N628), .Y(I228_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I158_un1_Y (.A(N555), .B(
        N483), .Y(I158_un1_Y));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I307_Y_0 (.A(off_div[17]), 
        .B(sum_39), .Y(ADD_32x32_fast_I307_Y_0));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I2_G0N (.A(sum_0_0), .B(
        \sum_adj[10]_net_1 ), .C(off_div[2]), .Y(N389));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I148_Y (.A(N536), .B(N533), 
        .C(N532), .Y(N597));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I48_Y (.A(off_div[21]), .B(
        off_div[22]), .C(sum_1_0), .Y(N494));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I260_un1_Y_0 (.A(N614), .B(
        N630), .Y(ADD_32x32_fast_I260_un1_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I33_Y (.A(off_div[29]), .B(
        off_div[30]), .C(sum_1_0), .Y(N479));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I268_un1_Y (.A(
        ADD_32x32_fast_I268_un1_Y_0), .B(N661), .Y(I268_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_3 (.A(N627), .B(N612), 
        .C(ADD_32x32_fast_I259_Y_2), .Y(ADD_32x32_fast_I259_Y_3));
    OR2B \off_div_RNIN351[5]  (.A(un5lto4), .B(off_div[5]), .Y(
        un1_off_divlt31));
    XNOR2 un1_nsum_adj_I_23 (.A(sum_8), .B(N_17), .Y(I_23_11));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I266_un1_Y_0 (.A(N642), .B(
        N626), .Y(ADD_32x32_fast_I266_un1_Y_0));
    XNOR2 un1_nsum_adj_I_28 (.A(sum_10), .B(N_15), .Y(I_28_3));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I67_Y (.A(off_div[12]), .B(
        \un1_sum_adj[12] ), .C(N423), .Y(N513));
    XNOR2 un1_nsum_adj_I_65 (.A(sum_22), .B(N_3), .Y(I_65_3));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I193_Y (.A(N582), .B(N590), 
        .Y(N648));
    OR2 \off_div_RNIRL7P[13]  (.A(off_div[13]), .B(off_div[14]), .Y(
        un5lto14_1));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I5_G0N (.A(\un1_sum_adj[5] )
        , .B(off_div[5]), .Y(N398));
    AND3 un1_nsum_adj_I_52 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[12] ), .Y(N_7));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I317_Y_0 (.A(off_div[27]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I317_Y_0));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y_1 (.A(I158_un1_Y), .B(
        N482), .C(I98_un1_Y), .Y(ADD_32x32_fast_I260_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I243_Y (.A(N644), .B(N659), 
        .C(N643), .Y(N784));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I296_Y_0 (.A(sum_2_0), .B(
        \sum_adj[14]_net_1 ), .C(off_div[6]), .Y(
        ADD_32x32_fast_I296_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I183_Y (.A(N572), .B(N580), 
        .Y(N638));
    NOR3 un1_nsum_adj_I_60 (.A(sum_19), .B(sum_18), .C(sum_20), .Y(
        \DWACT_FINC_E[15] ));
    MX2 \sum_adj_RNO[8]  (.A(sum_8), .B(I_23_11), .S(sum_0_0), .Y(
        \nsum_adj_5[8] ));
    XA1B \off_div_RNO[6]  (.A(N659), .B(ADD_32x32_fast_I296_Y_0), .C(
        \state[0]_net_1 ), .Y(\next_off_div[6] ));
    NOR3A \off_div_RNIA4KI1[26]  (.A(un1_off_divlto31_8), .B(
        off_div[26]), .C(off_div[27]), .Y(un1_off_divlto31_15));
    AO1C \state_RNI51T1I[1]  (.A(un5lt31), .B(next_off_div_2_sqmuxa_11)
        , .C(\state[1]_net_1 ), .Y(un1_state_2_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I124_Y (.A(N512), .B(N509), 
        .C(N508), .Y(N573));
    NOR2 un1_nsum_adj_I_21 (.A(sum_6), .B(sum_7), .Y(\DWACT_FINC_E[3] )
        );
    NOR2 \off_div_RNIPJ7P[13]  (.A(off_div[13]), .B(off_div[12]), .Y(
        un1_off_divlto31_2));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I201_Y (.A(N598), .B(N590), 
        .Y(N656));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I242_Y (.A(N642), .B(N657), 
        .C(N641), .Y(N781));
    DFN1E0C0 \off_div[1]  (.D(\next_off_div[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[1]));
    XA1 \off_div_RNO[8]  (.A(N802), .B(ADD_32x32_fast_I298_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[8] ));
    XNOR2 un1_nsum_adj_I_53 (.A(sum_18), .B(N_7), .Y(I_53_3));
    AND3 un1_nsum_adj_I_58 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[14] ), .Y(N_5));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I102_Y (.A(N490), .B(N486), 
        .Y(N551));
    MX2 \off_div_RNO[19]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[19] ), .S(\state_d[2] ), .Y(\next_off_div[19] ));
    DFN1E0C0 \off_div[10]  (.D(\next_off_div[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[10]));
    MX2 \off_div_RNO[10]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[10] ), .S(\state_d[2] ), .Y(\next_off_div[10] ));
    OR3 \off_div_RNII7FI1[11]  (.A(off_div[12]), .B(off_div[11]), .C(
        un5lto14_1), .Y(un5lto14_2));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I125_Y (.A(N509), .B(N513), 
        .Y(N574));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I263_Y_0 (.A(N561), .B(N554), 
        .C(N553), .Y(ADD_32x32_fast_I263_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I178_Y (.A(N575), .B(N568), 
        .C(N567), .Y(N633));
    DFN1E1C0 \sum_adj[12]  (.D(\nsum_adj_5[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[12]_net_1 ));
    XNOR2 un1_nsum_adj_I_49 (.A(sum_17), .B(N_8), .Y(I_49_3));
    MX2 \sum_adj_RNO[17]  (.A(sum_17), .B(I_49_3), .S(sum_0_0), .Y(
        \nsum_adj_5[17] ));
    NOR3A un1_nsum_adj_I_66 (.A(\DWACT_FINC_E[15] ), .B(sum_21), .C(
        sum_22), .Y(\DWACT_FINC_E[33] ));
    AND3 un1_nsum_adj_I_51 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[28] ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I297_Y (.A(\un1_sum_adj[7] ), 
        .B(off_div[7]), .C(N657), .Y(\un1_off_div_1[7] ));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I269_un1_Y (.A(N632), .B(
        N648), .C(N663), .Y(I269_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I136_Y (.A(N524), .B(N521), 
        .C(N520), .Y(N585));
    XA1B \off_div_RNO[16]  (.A(N779), .B(ADD_32x32_fast_I306_Y_0), .C(
        \state[0]_net_1 ), .Y(\next_off_div[16] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I35_Y (.A(off_div[28]), .B(
        off_div[29]), .C(sum_1_0), .Y(N481));
    MX2 \off_div_RNO[0]  (.A(next_off_div16), .B(\un1_off_div_1[0] ), 
        .S(\state_d_0[2] ), .Y(\next_off_div[0] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I199_Y (.A(N596), .B(N588), 
        .Y(N654));
    XA1 \off_div_RNO[23]  (.A(N765), .B(ADD_32x32_fast_I313_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[23] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I264_un1_Y_0 (.A(N622), .B(
        N638), .Y(ADD_32x32_fast_I264_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I87_Y (.A(N390), .B(N393), 
        .Y(N533));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I189_Y (.A(N586), .B(N578), 
        .Y(N644));
    MX2 \off_div_RNO[18]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[18] ), .S(\state_d[2] ), .Y(\next_off_div[18] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I38_Y (.A(off_div[26]), .B(
        off_div[27]), .C(sum_1_0), .Y(N484));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I187_Y (.A(N584), .B(N576), 
        .Y(N642));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I273_Y (.A(I273_un1_Y), .B(
        N639), .C(I240_un1_Y), .Y(N779));
    XA1 \off_div_RNO[25]  (.A(N761), .B(ADD_32x32_fast_I315_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[25] ));
    NOR3A \off_div_RNI2SJI1[24]  (.A(next_off_div_2_sqmuxa_3), .B(
        off_div[26]), .C(off_div[24]), .Y(next_off_div_2_sqmuxa_7));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I112_Y (.A(N500), .B(N496), 
        .Y(N561));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I14_G0N (.A(
        \un1_sum_adj[14] ), .B(off_div[14]), .Y(N425));
    DFN1E0C0 \off_div[12]  (.D(\next_off_div[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[12]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I271_Y_0 (.A(
        ADD_32x32_fast_I271_un1_Y_0), .B(N636), .C(N635), .Y(
        ADD_32x32_fast_I271_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I161_Y (.A(N550), .B(N558), 
        .Y(N616));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I103_Y (.A(N487), .B(N491), 
        .Y(N552));
    DFN1E0C0 \off_div[0]  (.D(\next_off_div[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[0]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I131_Y (.A(N519), .B(N515), 
        .Y(N580));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I120_Y (.A(N508), .B(N505), 
        .C(N504), .Y(N569));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I46_Y (.A(off_div[22]), .B(
        off_div[23]), .C(sum_1_0), .Y(N492));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I300_Y_0 (.A(off_div[10]), 
        .B(\sum_adj_RNIJIDD[18]_net_1 ), .Y(ADD_32x32_fast_I300_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I77_Y (.A(off_div[7]), .B(
        \un1_sum_adj[7] ), .C(N408), .Y(N523));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I44_Y (.A(off_div[23]), .B(
        off_div[24]), .C(sum_1_0), .Y(N490));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I260_Y_2 (.A(N614), .B(N629), 
        .C(ADD_32x32_fast_I260_Y_1), .Y(ADD_32x32_fast_I260_Y_2));
    AO1 \off_div_RNIUSQO8[31]  (.A(un1_off_divlto31_22), .B(
        un1_off_divlto31_21), .C(off_div[31]), .Y(next_off_div16));
    DFN1E1C0 \sum_adj[20]  (.D(\nsum_adj_5[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[20]_net_1 ));
    NOR3B \off_div_RNI4DKBD[30]  (.A(next_off_div_2_sqmuxa_9), .B(
        next_off_div_2_sqmuxa_8), .C(next_off_div16), .Y(
        next_off_div_2_sqmuxa_11));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I53_Y (.A(off_div[20]), .B(
        off_div[19]), .C(sum_2_0), .Y(N499));
    XOR2 \sum_adj_RNISORJ[12]  (.A(\sum_adj[12]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[4] ));
    MX2 \off_div_RNO[5]  (.A(next_off_div16), .B(\un1_off_div_1[5] ), 
        .S(\state_d_0[2] ), .Y(\next_off_div[5] ));
    XA1 \off_div_RNO[2]  (.A(N601), .B(ADD_32x32_fast_I292_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[2] ));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I6_G0N (.A(sum_0_0), .B(
        \sum_adj[14]_net_1 ), .C(off_div[6]), .Y(N401));
    NOR2 \state_RNIRC2F_2[1]  (.A(\state[1]_net_1 ), .B(
        \state[0]_net_1 ), .Y(pwm_rdy));
    NOR2 \off_div_RNI2V9P[25]  (.A(off_div[25]), .B(off_div[27]), .Y(
        next_off_div_2_sqmuxa_3));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I247_un1_Y (.A(N586), .B(
        N594), .C(N601), .Y(I247_un1_Y));
    XOR2 \sum_adj_RNITQSJ[22]  (.A(\sum_adj[22]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[14] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I151_Y (.A(N537), .B(
        \sum_adj_RNIH9EC[8]_net_1 ), .C(N536), .Y(N601));
    DFN1E0P0 \off_div[6]  (.D(\next_off_div[6] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[6]));
    DFN1E1C0 \sum_adj[17]  (.D(\nsum_adj_5[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[17]_net_1 ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I320_Y_0 (.A(off_div[30]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I320_Y_0));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I305_Y (.A(\un1_sum_adj[15] )
        , .B(off_div[15]), .C(N781), .Y(\un1_off_div_1[15] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I310_Y_0 (.A(off_div[20]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I310_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I270_Y_0 (.A(N649), .B(N634), 
        .C(N633), .Y(ADD_32x32_fast_I270_Y_0));
    AND3 un1_nsum_adj_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E[4] ));
    XOR2 \sum_adj_RNIURSJ[23]  (.A(\sum_adj[23]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[15] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I230_un1_Y (.A(N645), .B(
        N630), .Y(I230_un1_Y));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I52_Y (.A(off_div[19]), .B(
        off_div[20]), .C(sum_2_0), .Y(N498));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I204_Y (.A(I204_un1_Y), .B(
        N595), .Y(N661));
    NOR3A un1_nsum_adj_I_27 (.A(\DWACT_FINC_E[4] ), .B(sum_8), .C(
        sum_9), .Y(N_15));
    XOR2 \sum_adj_RNIJIDD[18]  (.A(\sum_adj[18]_net_1 ), .B(sum_2_0), 
        .Y(\sum_adj_RNIJIDD[18]_net_1 ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I263_un1_Y_0 (.A(N620), .B(
        N636), .Y(ADD_32x32_fast_I263_un1_Y_0));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y_0 (.A(N484), .B(
        I100_un1_Y), .Y(ADD_32x32_fast_I261_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I194_Y (.A(N591), .B(N584), 
        .C(N583), .Y(N649));
    NOR3A \off_div_RNIE3FI1[10]  (.A(un1_off_divlto31_2), .B(
        off_div[10]), .C(off_div[11]), .Y(un1_off_divlto31_12));
    NOR2 \off_div_RNIVSO[6]  (.A(off_div[6]), .B(off_div[7]), .Y(
        un1_off_divlto31_0));
    OA1 \off_div_RNI3DNE4[16]  (.A(off_div[16]), .B(un5lt16), .C(
        un5lto20_2), .Y(un5lt31));
    DFN1E0C0 \off_div[20]  (.D(\next_off_div[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[20]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I113_Y (.A(N501), .B(N497), 
        .Y(N562));
    NOR2A \state_RNIRC2F[1]  (.A(\state[1]_net_1 ), .B(
        \state[0]_net_1 ), .Y(\state_d_0[2] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I184_Y (.A(N581), .B(N574), 
        .C(N573), .Y(N639));
    NOR3C \off_div_RNIOG8J3[10]  (.A(un1_off_divlto31_13), .B(
        un1_off_divlto31_12), .C(un1_off_divlto31_17), .Y(
        un1_off_divlto31_21));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_0 (.A(off_div[28]), .B(
        off_div[29]), .C(sum_0_0), .Y(ADD_32x32_fast_I259_Y_0));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I294_Y_0 (.A(off_div[4]), .B(
        \un1_sum_adj[4] ), .Y(ADD_32x32_fast_I294_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I236_un1_Y (.A(N651), .B(
        N636), .Y(I236_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I10_G0N (.A(
        \sum_adj_RNIJIDD[18]_net_1 ), .B(off_div[10]), .Y(N413));
    XA1 \off_div_RNO[21]  (.A(N769), .B(ADD_32x32_fast_I311_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[21] ));
    DFN1E0C0 \off_div[18]  (.D(\next_off_div[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[18]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I262_un1_Y_0 (.A(N618), .B(
        N634), .Y(ADD_32x32_fast_I262_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I109_Y (.A(N497), .B(N493), 
        .Y(N558));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I146_Y (.A(N534), .B(N531), 
        .C(N530), .Y(N595));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I107_Y (.A(N491), .B(N495), 
        .Y(N556));
    AND3 un1_nsum_adj_I_54 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[9] ), .C(\DWACT_FINC_E[12] ), .Y(
        \DWACT_FINC_E[13] ));
    AND3 un1_nsum_adj_I_69 (.A(\DWACT_FINC_E[29] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[33] ), .Y(N_2));
    NOR2 \off_div_RNIVR9P[24]  (.A(off_div[24]), .B(off_div[25]), .Y(
        un1_off_divlto31_10));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I195_Y (.A(N592), .B(N584), 
        .Y(N650));
    NOR2 un1_nsum_adj_I_57 (.A(sum_18), .B(sum_19), .Y(
        \DWACT_FINC_E[14] ));
    XOR2 \sum_adj_RNIH9EC[8]  (.A(\sum_adj[8]_net_1 ), .B(sum_39), .Y(
        \sum_adj_RNIH9EC[8]_net_1 ));
    NOR2 \off_div_RNI74AP[28]  (.A(off_div[28]), .B(off_div[29]), .Y(
        un1_off_divlto31_8));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I63_Y (.A(N429), .B(N426), 
        .Y(N509));
    NOR2A un1_nsum_adj_I_25 (.A(\DWACT_FINC_E[4] ), .B(sum_8), .Y(N_16)
        );
    DFN1E0C0 \off_div[22]  (.D(\next_off_div[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[22]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I185_Y (.A(N574), .B(N582), 
        .Y(N640));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I90_Y (.A(N383), .B(N387), .C(
        N386), .Y(N536));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I55_Y (.A(off_div[19]), .B(
        off_div[18]), .C(sum_2_0), .Y(N501));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I49_Y (.A(off_div[22]), .B(
        off_div[21]), .C(sum_1_0), .Y(N495));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I259_Y_2 (.A(N553), .B(N546), 
        .C(ADD_32x32_fast_I259_Y_1), .Y(ADD_32x32_fast_I259_Y_2));
    XA1 \off_div_RNO[12]  (.A(N790), .B(ADD_32x32_fast_I302_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[12] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I62_Y (.A(N425), .B(N429), .C(
        N428), .Y(N508));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y (.A(
        ADD_32x32_fast_I261_un1_Y_0), .B(N790), .C(
        ADD_32x32_fast_I261_Y_2), .Y(N755));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I141_Y (.A(N529), .B(N525), 
        .Y(N590));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I36_Y (.A(off_div[27]), .B(
        off_div[28]), .C(sum_1_0), .Y(N482));
    NOR3C \off_div_RNIHNOJ1[5]  (.A(un1_off_divlto31_10), .B(
        un1_off_divlto31_9), .C(un1_off_divlt31), .Y(
        un1_off_divlto31_20));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I58_Y (.A(off_div[16]), .B(
        off_div[17]), .C(sum_2_0), .Y(N504));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I292_Y_0 (.A(sum_2_0), .B(
        \sum_adj[10]_net_1 ), .C(off_div[2]), .Y(
        ADD_32x32_fast_I292_Y_0));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I91_Y (.A(sum_0_0), .B(
        off_div[0]), .C(N387), .Y(N537));
    DFN1E0C0 \off_div[17]  (.D(\next_off_div[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[17]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I119_Y (.A(N503), .B(N507), 
        .Y(N568));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I190_Y (.A(I190_un1_Y), .B(
        N579), .Y(N645));
    MX2 \sum_adj_RNO[23]  (.A(sum_23), .B(I_70_3), .S(sum_1_0), .Y(
        \nsum_adj_5[23] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I117_Y (.A(N501), .B(N505), 
        .Y(N566));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I132_Y (.A(N520), .B(N517), 
        .C(N516), .Y(N581));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I180_Y (.A(N577), .B(N570), 
        .C(N569), .Y(N635));
    NOR3B un1_nsum_adj_I_55 (.A(\DWACT_FINC_E[13] ), .B(
        \DWACT_FINC_E[28] ), .C(sum_18), .Y(N_6));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I128_Y (.A(N516), .B(N513), 
        .C(N512), .Y(N577));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I104_Y (.A(N492), .B(
        I100_un1_Y), .Y(N553));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I240_un1_Y (.A(N655), .B(
        N640), .Y(I240_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I15_G0N (.A(
        \un1_sum_adj[15] ), .B(off_div[15]), .Y(N428));
    XOR2 \sum_adj_RNIVRRJ[15]  (.A(\sum_adj[15]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[7] ));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I273_un1_Y (.A(N656), .B(
        \sum_adj_RNIH9EC[8]_net_1 ), .C(N640), .Y(I273_un1_Y));
    NOR3 un1_nsum_adj_I_50 (.A(sum_17), .B(sum_16), .C(sum_15), .Y(
        \DWACT_FINC_E[12] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I295_Y_0 (.A(off_div[5]), .B(
        \un1_sum_adj[5] ), .Y(ADD_32x32_fast_I295_Y_0));
    NOR2 \off_div_RNIRN9P[22]  (.A(off_div[22]), .B(off_div[23]), .Y(
        un1_off_divlto31_9));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I176_Y (.A(N573), .B(N566), 
        .C(N565), .Y(N631));
    XNOR2 un1_nsum_adj_I_26 (.A(sum_9), .B(N_16), .Y(I_26_3));
    DFN1E0C0 \off_div[28]  (.D(\next_off_div[28] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[28]));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I83_Y (.A(off_div[5]), .B(
        \un1_sum_adj[5] ), .C(N396), .Y(N529));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I65_Y (.A(N426), .B(N423), 
        .Y(N511));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I246_un1_Y (.A(N650), .B(
        N599), .Y(I246_un1_Y));
    DFN1C0 \state[1]  (.D(N_311_i), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \state[1]_net_1 ));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I15_P0N (.A(\un1_sum_adj[15] )
        , .B(off_div[15]), .Y(N429));
    XA1B \off_div_RNO[31]  (.A(N749), .B(ADD_32x32_fast_I321_Y_0), .C(
        \state[0]_net_1 ), .Y(\next_off_div[31] ));
    XA1 \off_div_RNO[14]  (.A(N784), .B(ADD_32x32_fast_I304_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[14] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I105_Y (.A(N489), .B(N493), 
        .Y(N554));
    NOR2A \state_RNIRC2F_1[1]  (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(state_176_d));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I163_Y (.A(N552), .B(N560), 
        .Y(N618));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I133_Y (.A(N517), .B(N521), 
        .Y(N582));
    NOR2 \off_div_RNI508P[18]  (.A(off_div[18]), .B(off_div[19]), .Y(
        un1_off_divlto31_4));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I190_un1_Y (.A(N587), .B(
        N580), .Y(I190_un1_Y));
    XOR2 \sum_adj_RNI0TRJ[16]  (.A(\sum_adj[16]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[8] ));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I68_Y (.A(N416), .B(
        off_div[12]), .C(\un1_sum_adj[12] ), .Y(N514));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I114_Y (.A(N502), .B(N498), 
        .Y(N563));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I261_un1_Y_0 (.A(N616), .B(
        N632), .Y(ADD_32x32_fast_I261_un1_Y_0));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I82_Y (.A(N395), .B(
        off_div[5]), .C(\un1_sum_adj[5] ), .Y(N528));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I171_Y (.A(N560), .B(N568), 
        .Y(N626));
    NOR3 un1_nsum_adj_I_18 (.A(sum_4), .B(sum_3), .C(sum_5), .Y(
        \DWACT_FINC_E[2] ));
    MX2 \sum_adj_RNO[14]  (.A(sum_14), .B(I_40_3), .S(sum_0_0), .Y(
        \nsum_adj_5[14] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I40_Y (.A(off_div[26]), .B(
        off_div[25]), .C(sum_1_0), .Y(N486));
    DFN1E1C0 \sum_adj[8]  (.D(\nsum_adj_5[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[8]_net_1 ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I204_un1_Y (.A(N596), .B(
        N538), .Y(I204_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I12_G0N (.A(
        \un1_sum_adj[12] ), .B(off_div[12]), .Y(N419));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I11_P0N (.A(sum_1_0), .B(
        \sum_adj[19]_net_1 ), .C(off_div[11]), .Y(N417));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I73_Y (.A(off_div[9]), .B(
        \un1_sum_adj[9] ), .C(N414), .Y(N519));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I266_Y_0 (.A(N641), .B(N626), 
        .C(N625), .Y(ADD_32x32_fast_I266_Y_0));
    OR2 \off_div_RNIPMO[3]  (.A(off_div[4]), .B(off_div[3]), .Y(
        un5lto4));
    XNOR2 un1_nsum_adj_I_56 (.A(sum_19), .B(N_6), .Y(I_56_3));
    OA1B \state_RNO[0]  (.A(\state[1]_net_1 ), .B(pwm_enable), .C(
        \state[0]_net_1 ), .Y(\state_ns[0] ));
    DFN1E0C0 \off_div[2]  (.D(\next_off_div[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[2]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I39_Y (.A(off_div[27]), .B(
        off_div[26]), .C(sum_1_0), .Y(N485));
    DFN1E0C0 \off_div[27]  (.D(\next_off_div[27] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[27]));
    MX2 \sum_adj_RNO[18]  (.A(sum_18), .B(I_53_3), .S(sum_0_0), .Y(
        \nsum_adj_5[18] ));
    DFN1E1C0 \sum_adj[15]  (.D(\nsum_adj_5[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[15]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I41_Y (.A(off_div[25]), .B(
        off_div[26]), .C(sum_1_0), .Y(N487));
    XNOR2 un1_nsum_adj_I_32 (.A(sum_11), .B(N_14), .Y(I_32_3));
    XOR2 \sum_adj_RNI1URJ[17]  (.A(\sum_adj[17]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[9] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I264_Y (.A(
        ADD_32x32_fast_I264_un1_Y_0), .B(N799), .C(
        ADD_32x32_fast_I264_Y_1), .Y(N761));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I72_Y (.A(N410), .B(N414), .C(
        N413), .Y(N518));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I295_Y (.A(
        ADD_32x32_fast_I295_Y_0), .B(N661), .Y(\un1_off_div_1[5] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I262_un1_Y (.A(
        ADD_32x32_fast_I262_un1_Y_0), .B(N793), .Y(I262_un1_Y));
    XA1 \off_div_RNO[29]  (.A(N753), .B(ADD_32x32_fast_I319_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[29] ));
    DFN1E0C0 \off_div[14]  (.D(\next_off_div[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[14]));
    DFN1E1C0 \sum_adj[10]  (.D(\nsum_adj_5[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[10]_net_1 ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I302_Y_0 (.A(off_div[12]), 
        .B(\un1_sum_adj[12] ), .Y(ADD_32x32_fast_I302_Y_0));
    MX2 \off_div_RNO[20]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[20] ), .S(\state_d[2] ), .Y(\next_off_div[20] ));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I300_Y (.A(
        ADD_32x32_fast_I300_Y_0), .B(N796), .Y(\un1_off_div_1[10] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I115_Y (.A(N499), .B(N503), 
        .Y(N564));
    XOR2 \sum_adj_RNITPRJ[13]  (.A(\sum_adj[13]_net_1 ), .B(sum_39), 
        .Y(\un1_sum_adj[5] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I258_un1_Y_0 (.A(N610), .B(
        N626), .Y(ADD_32x32_fast_I258_un1_Y_0));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I142_Y (.A(N530), .B(N527), 
        .C(N526), .Y(N591));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I56_Y (.A(off_div[17]), .B(
        off_div[18]), .C(sum_2_0), .Y(N502));
    XA1 \off_div_RNO[26]  (.A(N759), .B(ADD_32x32_fast_I316_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[26] ));
    NOR3C \off_div_RNIMA853[24]  (.A(un1_off_divlto31_9), .B(
        next_off_div_2_sqmuxa_0), .C(next_off_div_2_sqmuxa_7), .Y(
        next_off_div_2_sqmuxa_9));
    MX2 \sum_adj_RNO[13]  (.A(sum_13), .B(I_37_3), .S(sum_0_0), .Y(
        \nsum_adj_5[13] ));
    DFN1E1C0 \sum_adj[19]  (.D(\nsum_adj_5[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[19]_net_1 ));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I267_un1_Y (.A(N628), .B(
        N644), .C(N659), .Y(I267_un1_Y));
    XOR2 \sum_adj_RNIIAEC[9]  (.A(\sum_adj[9]_net_1 ), .B(sum_39), .Y(
        \un1_sum_adj[1] ));
    MX2 \off_div_RNO[17]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[17] ), .S(\state_d[2] ), .Y(\next_off_div[17] ));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I54_Y (.A(off_div[18]), .B(
        off_div[19]), .C(sum_2_0), .Y(N500));
    OR3 un1_off_div_1_0_0_ADD_32x32_fast_I267_Y (.A(I228_un1_Y), .B(
        N627), .C(I267_un1_Y), .Y(N767));
    DFN1E0C0 \off_div[4]  (.D(\next_off_div[4] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[4]));
    NOR3 un1_nsum_adj_I_33 (.A(sum_10), .B(sum_9), .C(sum_11), .Y(
        \DWACT_FINC_E[7] ));
    NOR2 un1_nsum_adj_I_38 (.A(sum_12), .B(sum_13), .Y(
        \DWACT_FINC_E[8] ));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I303_Y_0 (.A(sum_1_0), .B(
        \sum_adj[21]_net_1 ), .C(off_div[13]), .Y(
        ADD_32x32_fast_I303_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I169_Y (.A(N566), .B(N558), 
        .Y(N624));
    DFN1E0C0 \off_div[19]  (.D(\next_off_div[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[19]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I85_Y (.A(N396), .B(N393), 
        .Y(N531));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I312_Y_0 (.A(off_div[22]), 
        .B(sum_39), .Y(ADD_32x32_fast_I312_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I268_un1_Y_0 (.A(N646), .B(
        N630), .Y(ADD_32x32_fast_I268_un1_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I139_Y (.A(N527), .B(N523), 
        .Y(N588));
    XA1 \off_div_RNO[28]  (.A(N755), .B(ADD_32x32_fast_I318_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[28] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I167_Y (.A(N564), .B(N556), 
        .Y(N622));
    NOR3A \off_div_RNISJHI1[20]  (.A(un1_off_divlto31_4), .B(
        off_div[20]), .C(off_div[21]), .Y(un1_off_divlto31_13));
    DFN1E0C0 \off_div[16]  (.D(\next_off_div[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[16]));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I8_P0N (.A(\un1_sum_adj[8] ), 
        .B(off_div[8]), .Y(N408));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I198_Y (.A(N595), .B(N588), 
        .C(N587), .Y(N653));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I137_Y (.A(N521), .B(N525), 
        .Y(N586));
    DFN1E0C0 \off_div[8]  (.D(\next_off_div[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[8]));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I97_Y (.A(N485), .B(N481), 
        .Y(N546));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I188_Y (.A(N585), .B(N578), 
        .C(N577), .Y(N643));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I16_P0N (.A(off_div[16]), .B(
        sum_39), .Y(N432));
    OR2 un1_off_div_1_0_0_ADD_32x32_fast_I110_Y (.A(N498), .B(N494), 
        .Y(I162_un1_Y));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I88_Y (.A(N386), .B(N390), .C(
        N389), .Y(N534));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_0 (.A(off_div[30]), .B(
        off_div[29]), .C(sum_2_0), .Y(ADD_32x32_fast_I258_Y_0));
    NOR3 un1_nsum_adj_I_29 (.A(sum_7), .B(sum_6), .C(sum_8), .Y(
        \DWACT_FINC_E[5] ));
    NOR3A \off_div_RNIUJFI1[16]  (.A(un1_off_divlto31_6), .B(
        off_div[16]), .C(off_div[17]), .Y(un1_off_divlto31_14));
    AX1D un1_off_div_1_0_0_ADD_32x32_fast_I310_Y (.A(I269_un1_Y), .B(
        ADD_32x32_fast_I269_Y_0), .C(ADD_32x32_fast_I310_Y_0), .Y(
        \un1_off_div_1[20] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y_2 (.A(N616), .B(N631), 
        .C(ADD_32x32_fast_I261_Y_1), .Y(ADD_32x32_fast_I261_Y_2));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I159_Y (.A(N483), .B(N487), 
        .C(N556), .Y(N614));
    NOR3A un1_nsum_adj_I_31 (.A(\DWACT_FINC_E[6] ), .B(sum_9), .C(
        sum_10), .Y(N_14));
    OA1 \off_div_RNIINIF2[15]  (.A(un5lt14), .B(un5lto14_2), .C(
        off_div[15]), .Y(un5lt16));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I313_Y_0 (.A(off_div[23]), 
        .B(sum_2_0), .Y(ADD_32x32_fast_I313_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I157_Y (.A(N546), .B(N554), 
        .Y(N612));
    OA1 un1_off_div_1_0_0_ADD_32x32_fast_I75_Y (.A(off_div[9]), .B(
        \un1_sum_adj[9] ), .C(N408), .Y(N521));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I293_Y (.A(
        ADD_32x32_fast_I293_Y_0), .B(N599), .Y(\un1_off_div_1[3] ));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I143_Y (.A(N527), .B(N531), 
        .Y(N592));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I259_un1_Y_0 (.A(N612), .B(
        N628), .Y(ADD_32x32_fast_I259_un1_Y_0));
    DFN1E0P0 \off_div[3]  (.D(\next_off_div[3] ), .CLK(clk_c), .PRE(
        n_rst_c), .E(un1_state_2_0), .Q(off_div[3]));
    XOR3 un1_off_div_1_0_0_ADD_32x32_fast_I290_Y (.A(sum_1_0), .B(
        off_div[0]), .C(\sum_adj_RNIH9EC[8]_net_1 ), .Y(
        \un1_off_div_1[0] ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_1 (.A(N479), .B(N482), 
        .C(ADD_32x32_fast_I258_Y_0), .Y(ADD_32x32_fast_I258_Y_1));
    MX2 \off_div_RNO[7]  (.A(next_off_div_1_sqmuxa), .B(
        \un1_off_div_1[7] ), .S(\state_d_0[2] ), .Y(\next_off_div[7] ));
    MAJ3 un1_off_div_1_0_0_ADD_32x32_fast_I78_Y (.A(N401), .B(
        off_div[7]), .C(\un1_sum_adj[7] ), .Y(N524));
    NOR3A \off_div_RNIEP7E[30]  (.A(un1_off_divlto31_0), .B(
        off_div[30]), .C(un5lto9), .Y(un1_off_divlto31_17));
    DFN1E1C0 \sum_adj[21]  (.D(\nsum_adj_5[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[21]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I258_Y_3 (.A(N625), .B(N610), 
        .C(ADD_32x32_fast_I258_Y_2), .Y(ADD_32x32_fast_I258_Y_3));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I66_Y (.A(N419), .B(N423), .C(
        N422), .Y(N512));
    NOR3C un1_off_div_1_0_0_ADD_32x32_fast_I270_un1_Y (.A(N634), .B(
        N650), .C(N599), .Y(I270_un1_Y));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I8_G0N (.A(\un1_sum_adj[8] )
        , .B(off_div[8]), .Y(N407));
    XOR2 un1_off_div_1_0_0_ADD_32x32_fast_I299_Y_0 (.A(off_div[9]), .B(
        \un1_sum_adj[9] ), .Y(ADD_32x32_fast_I299_Y_0));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I1_G0N (.A(\un1_sum_adj[1] )
        , .B(off_div[1]), .Y(N386));
    XA1 \off_div_RNO[4]  (.A(N663), .B(ADD_32x32_fast_I294_Y_0), .C(
        \state_d_0[2] ), .Y(\next_off_div[4] ));
    DFN1E0C0 \off_div[24]  (.D(\next_off_div[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_RNI51T1I_0[1]_net_1 ), .Q(off_div[24]));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I64_Y (.A(N422), .B(N426), .C(
        N425), .Y(N510));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I205_Y (.A(N598), .B(
        \sum_adj_RNIH9EC[8]_net_1 ), .C(N597), .Y(N663));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I172_Y (.A(N569), .B(N562), 
        .C(N561), .Y(N627));
    XNOR2 un1_nsum_adj_I_59 (.A(sum_20), .B(N_5), .Y(I_59_3));
    OR2 \off_div_RNI31P[8]  (.A(off_div[8]), .B(off_div[9]), .Y(
        un5lto9));
    XA1 un1_off_div_1_0_0_ADD_32x32_fast_I3_G0N (.A(sum_1_0), .B(
        \sum_adj[11]_net_1 ), .C(off_div[3]), .Y(N392));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I134_Y (.A(N522), .B(N519), 
        .C(N518), .Y(N583));
    AND3 un1_nsum_adj_I_42 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[9] ), .Y(N_10));
    DFN1E1C0 \sum_adj[16]  (.D(\nsum_adj_5[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(state_176_d), .Q(\sum_adj[16]_net_1 ));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I244_Y (.A(N646), .B(N661), 
        .C(N645), .Y(N787));
    NOR2B un1_off_div_1_0_0_ADD_32x32_fast_I238_un1_Y (.A(N653), .B(
        N638), .Y(I238_un1_Y));
    MX2 \sum_adj_RNO[19]  (.A(sum_19), .B(I_56_3), .S(sum_0_0), .Y(
        \nsum_adj_5[19] ));
    XO1 un1_off_div_1_0_0_ADD_32x32_fast_I6_P0N (.A(sum_0_0), .B(
        \sum_adj[14]_net_1 ), .C(off_div[6]), .Y(N402));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I261_Y_1 (.A(N557), .B(N550), 
        .C(ADD_32x32_fast_I261_Y_0), .Y(ADD_32x32_fast_I261_Y_1));
    AO1 un1_off_div_1_0_0_ADD_32x32_fast_I126_Y (.A(N514), .B(N511), 
        .C(N510), .Y(N575));
    XA1 \off_div_RNO[30]  (.A(N751), .B(ADD_32x32_fast_I320_Y_0), .C(
        \state_d[2] ), .Y(\next_off_div[30] ));
    
endmodule


module integral_calc_13s_4_3(
       avg_old,
       avg_new,
       average,
       LED_15,
       LED_15_i_0,
       calc_avg,
       N_46_1,
       n_rst_c,
       clk_c
    );
input  [11:0] avg_old;
input  [11:0] avg_new;
output [6:2] average;
output [7:0] LED_15;
output LED_15_i_0;
input  calc_avg;
output N_46_1;
input  n_rst_c;
input  clk_c;

    wire \state_1[0]_net_1 , \state_1_RNIDTBQ[0]_net_1 , 
        \state_0[0]_net_1 , N637, N521, I188_un1_Y, N643, N525, 
        I190_un1_Y, N649, N529, I192_un1_Y, N640, N523, I189_un1_Y, 
        \un1_integ[14] , ADD_26x26_fast_I244_Y_0, \un1_integ[13] , 
        ADD_26x26_fast_I243_Y_0, \un1_integ[15] , 
        ADD_26x26_fast_I245_Y_0, \integ[15]_net_1 , \state[0]_net_1 , 
        ADD_26x26_fast_I241_Y_0, \un1_next_int[11] , \un1_integ[11] , 
        ADD_26x26_fast_I253_Y_0, \integ[23]_net_1 , 
        ADD_26x26_fast_I254_Y_0, \integ[24]_net_1 , 
        ADD_26x26_fast_I255_Y_0, \integ[25]_net_1 , 
        ADD_26x26_fast_I206_Y_2, N506, ADD_26x26_fast_I206_Y_1, N402, 
        N398, N459, ADD_26x26_fast_I252_Y_0, \integ[22]_net_1 , 
        ADD_26x26_fast_I204_Y_3, N502, N517, ADD_26x26_fast_I204_Y_2, 
        ADD_26x26_fast_I204_Y_0, N455, ADD_26x26_fast_I205_Y_3, N504, 
        N519, ADD_26x26_fast_I205_Y_2, N400, ADD_26x26_fast_I205_Y_0, 
        N457, ADD_26x26_fast_I251_Y_0, \integ[21]_net_1 , 
        ADD_26x26_fast_I250_Y_0, \integ[20]_net_1 , 
        ADD_26x26_fast_I237_Y_0, \un1_next_int[7] , 
        ADD_26x26_fast_I249_Y_0, \integ[19]_net_1 , 
        ADD_26x26_fast_I207_Y_2, N508, ADD_26x26_fast_I207_Y_1, N404, 
        N461, ADD_26x26_fast_I248_Y_0, \integ[18]_net_1 , 
        ADD_26x26_fast_I209_Y_1, ADD_26x26_fast_I209_un1_Y_0, N543, 
        ADD_26x26_fast_I209_Y_0, N465, N458, ADD_26x26_fast_I208_Y_1, 
        ADD_26x26_fast_I208_un1_Y_0, N541, ADD_26x26_fast_I208_Y_0, 
        N463, ADD_26x26_fast_I239_Y_0, \un18_next_int_m[9] , 
        \inf_abs0_m[9] , ADD_26x26_fast_I238_Y_0, \inf_abs0_m[8] , 
        \un18_next_int_m[8] , ADD_26x26_fast_I210_Y_1, 
        ADD_26x26_fast_I210_un1_Y_0, N491, ADD_26x26_fast_I210_Y_0, 
        N467, N460, ADD_26x26_fast_I204_un1_Y_0, N472, N464, 
        ADD_26x26_fast_I205_un1_Y_0, N520, ADD_26x26_fast_I240_Y_0, 
        \un1_next_int[10] , ADD_26x26_fast_I211_Y_1, 
        ADD_26x26_fast_I211_un1_Y_0, N516, ADD_26x26_fast_I211_Y_0, 
        N469, N462, ADD_26x26_fast_I213_Y_0, 
        ADD_26x26_fast_I213_un1_Y_0, ADD_26x26_fast_I207_un1_Y_0, N478, 
        N470, ADD_26x26_fast_I234_Y_0, \un1_next_int[4] , 
        ADD_26x26_fast_I235_Y_0, \un18_next_int_m[5] , \inf_abs0_m[5] , 
        N512, N528, N510, N526, ADD_26x26_fast_I233_Y_0, 
        \un18_next_int_m[3] , \inf_abs0_m[3] , N476, N484, N514, 
        ADD_26x26_fast_I212_un1_Y_0, N480, N488, N442, N482, N490, 
        \un1_next_int[0] , N486, N493, ADD_26x26_fast_I232_Y_0, 
        \un1_next_int[2] , ADD_26x26_fast_I127_Y_1, 
        ADD_26x26_fast_I127_Y_0, N401, ADD_26x26_fast_I125_Y_0, 
        ADD_26x26_fast_I230_Y_2, \state[1]_net_1 , \integ[0]_net_1 , 
        \un1_integ[18] , I182_un1_Y, \un1_integ[20] , I178_un1_Y, 
        \un1_integ[19] , I180_un1_Y, \un1_integ[24] , I205_un1_Y, 
        \un1_integ[23] , I206_un1_Y, N522, N537, N399, N403, N535, 
        I195_un1_Y, ADD_26x26_fast_I238_Y, N633, I212_un1_Y, 
        I184_un1_Y, \un1_integ[17] , \integ[17]_net_1 , 
        \un1_integ[25] , I204_un1_Y, ADD_26x26_fast_I236_Y, 
        \un1_next_int[6] , N539, ADD_26x26_fast_I242_Y, N646, 
        \un1_integ[16] , \integ[16]_net_1 , N635, 
        ADD_26x26_fast_I233_Y_0_0, ADD_26x26_fast_I237_Y, 
        \un1_integ[21] , I176_un1_Y, ADD_26x26_fast_I232_Y_0_0, 
        ADD_26x26_fast_I240_Y, N531, I193_un1_Y, \un1_integ[22] , 
        I207_un1_Y, ADD_26x26_fast_I239_Y, N533, I194_un1_Y, 
        ADD_26x26_fast_I235_Y, ADD_26x26_fast_I234_Y_0_0, 
        ADD_26x26_fast_I231_Y_0, \un1_next_int[1] , \integ[1]_net_1 , 
        N405, N456, N474, N489, N481, I163_un1_Y, N527, N487, N479, 
        N430, N427, N426, N338, N342, N341, N339, N431, N333, N439, 
        N435, N327, N321, N324, I150_un1_Y, N473, N424, N421, N420, 
        N425, N345, N477, N417, N416, N429, N466, N413, N363, N366, 
        N415, N423, N348, N471, N414, N410, N440, N437, N436, N323, 
        N326, N441, N318, N433, N432, N428, N335, N332, N317, N483, 
        N434, N438, I120_un1_Y, I148_un1_Y, I162_un1_Y, N418, N407, 
        N320, N329, N347, N344, N485, I121_un1_Y, \un18_next_int_m[0] , 
        \inf_abs0_m[4] , \un18_next_int_m[4] , \inf_abs0_m[7] , 
        \un18_next_int_m[7] , \inf_abs0_m[10] , \un18_next_int_m[10] , 
        \inf_abs0_m[11] , \un18_next_int_m[11] , \inf_abs0_m[1] , 
        \un18_next_int_m[1] , \inf_abs0_m[2] , \un18_next_int_m[2] , 
        \inf_abs0_m[6] , \un18_next_int_m[6] , \state_RNO_7[1] , N409, 
        N362, N412, N359, N422, N350, N354, N353, N360, N357, N351, 
        N356, I152_un1_Y, N475, N468, N419, N408, N406, GND, VCC;
    
    AO1 un1_integ_0_0_ADD_26x26_fast_I56_Y (.A(N341), .B(N345), .C(
        N344), .Y(N424));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I148_un1_Y (.A(N479), .B(N472), 
        .Y(I148_un1_Y));
    OR2A un1_integ_0_0_ADD_26x26_fast_I15_P0N (.A(\state[0]_net_1 ), 
        .B(\integ[15]_net_1 ), .Y(N363));
    DFN1C0 \state[0]  (.D(\state_1_RNIDTBQ[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state[0]_net_1 ));
    DFN1E0C0 \integ[13]  (.D(\un1_integ[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(LED_15[6]));
    DFN1E0C0 \integ[24]  (.D(\un1_integ[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(\integ[24]_net_1 ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I245_Y_0 (.A(\integ[15]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I245_Y_0));
    OA1 un1_integ_0_0_ADD_26x26_fast_I61_Y (.A(average[6]), .B(
        \un1_next_int[6] ), .C(N339), .Y(N429));
    OR2 un1_integ_0_0_ADD_26x26_fast_I7_P0N (.A(\un1_next_int[7] ), .B(
        LED_15[0]), .Y(N339));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I248_Y_0 (.A(\integ[18]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I248_Y_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I41_Y (.A(\integ[17]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_1[0]_net_1 ), .Y(N409));
    OA1 un1_integ_0_0_ADD_26x26_fast_I204_un1_Y (.A(N533), .B(
        I194_un1_Y), .C(ADD_26x26_fast_I204_un1_Y_0), .Y(I204_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I86_Y (.A(N404), .B(N408), .Y(
        N457));
    AO1 un1_integ_0_0_ADD_26x26_fast_I98_Y (.A(N420), .B(N417), .C(
        N416), .Y(N469));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I176_un1_Y (.A(N510), .B(N525), 
        .Y(I176_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I205_un1_Y_0 (.A(N504), .B(N520)
        , .Y(ADD_26x26_fast_I205_un1_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I150_un1_Y (.A(N481), .B(N474), 
        .Y(I150_un1_Y));
    NOR2A un1_integ_0_0_ADD_26x26_fast_I14_G0N (.A(LED_15[7]), .B(
        \state[0]_net_1 ), .Y(N359));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I51_Y (.A(N354), .B(N351), .Y(
        N419));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I230_Y (.A(\state[1]_net_1 ), .B(
        \integ[0]_net_1 ), .C(\un1_next_int[0] ), .Y(
        ADD_26x26_fast_I230_Y_2));
    NOR2A \state_RNIAGJR[1]  (.A(\state[1]_net_1 ), .B(avg_old[11]), 
        .Y(\un18_next_int_m[11] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I253_Y (.A(I206_un1_Y), .B(
        ADD_26x26_fast_I206_Y_2), .C(ADD_26x26_fast_I253_Y_0), .Y(
        \un1_integ[23] ));
    DFN1E0C0 \integ[21]  (.D(\un1_integ[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(\integ[21]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I190_un1_Y (.A(N526), .B(N541), 
        .Y(I190_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I146_Y (.A(N477), .B(N470), .C(
        N469), .Y(N523));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I210_un1_Y_0 (.A(N476), .B(N484)
        , .C(N514), .Y(ADD_26x26_fast_I210_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I142_Y (.A(N473), .B(N466), .C(
        N465), .Y(N519));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I244_Y_0 (.A(LED_15[7]), .B(
        \state_1[0]_net_1 ), .Y(ADD_26x26_fast_I244_Y_0));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I231_Y (.A(\un1_next_int[1] ), 
        .B(\integ[1]_net_1 ), .C(N442), .Y(ADD_26x26_fast_I231_Y_0));
    DFN1E0C0 \integ[15]  (.D(\un1_integ[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(\integ[15]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I103_Y (.A(N421), .B(N425), .Y(
        N474));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I125_Y (.A(N399), .B(
        ADD_26x26_fast_I125_Y_0), .C(N456), .Y(N502));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_1 (.A(
        ADD_26x26_fast_I209_un1_Y_0), .B(N543), .C(
        ADD_26x26_fast_I209_Y_0), .Y(ADD_26x26_fast_I209_Y_1));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I97_Y (.A(N415), .B(N419), .Y(
        N468));
    AO1 un1_integ_0_0_ADD_26x26_fast_I94_Y (.A(N416), .B(N413), .C(
        N412), .Y(N465));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I151_Y (.A(N482), .B(N474), .Y(
        N528));
    AO1 un1_integ_0_0_ADD_26x26_fast_I74_Y (.A(N318), .B(
        \un1_next_int[0] ), .C(N317), .Y(N442));
    AX1D un1_integ_0_0_ADD_26x26_fast_I238_Y (.A(N535), .B(I195_un1_Y), 
        .C(ADD_26x26_fast_I238_Y_0), .Y(ADD_26x26_fast_I238_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I121_Y (.A(I121_un1_Y), .B(N440), 
        .Y(N493));
    OR2 \state_RNIJ87F1[0]  (.A(\inf_abs0_m[4] ), .B(
        \un18_next_int_m[4] ), .Y(\un1_next_int[4] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I190_Y (.A(N525), .B(I190_un1_Y), 
        .Y(N643));
    OR3 un1_integ_0_0_ADD_26x26_fast_I5_P0N (.A(\un18_next_int_m[5] ), 
        .B(\inf_abs0_m[5] ), .C(average[5]), .Y(N333));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I246_Y (.A(\state_0[0]_net_1 ), 
        .B(\integ[16]_net_1 ), .C(N635), .Y(\un1_integ[16] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I252_Y_0 (.A(\integ[22]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I252_Y_0));
    DFN1C0 \state_1[0]  (.D(\state_1_RNIDTBQ[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_1[0]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I39_Y (.A(\integ[17]_net_1 ), .B(
        \integ[18]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N407));
    OA1B un1_integ_0_0_ADD_26x26_fast_I32_Y (.A(\integ[20]_net_1 ), .B(
        \integ[21]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N400));
    AO1 un1_integ_0_0_ADD_26x26_fast_I213_Y (.A(N535), .B(N520), .C(
        ADD_26x26_fast_I213_Y_0), .Y(N635));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I194_un1_Y (.A(N480), .B(N488), 
        .C(N442), .Y(I194_un1_Y));
    AO1B un1_integ_0_0_ADD_26x26_fast_I125_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\integ[24]_net_1 ), .C(\state_0[0]_net_1 ), .Y(
        ADD_26x26_fast_I125_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I100_Y (.A(N422), .B(N419), .C(
        N418), .Y(N471));
    OR2 un1_integ_0_0_ADD_26x26_fast_I12_P0N (.A(LED_15[5]), .B(
        \state[1]_net_1 ), .Y(N354));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I10_G0N (.A(\un1_next_int[10] ), 
        .B(LED_15[3]), .Y(N347));
    NOR2B \state_RNIK87N[0]  (.A(avg_new[1]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[1] ));
    OR2 \state_1_RNIVSNB1[0]  (.A(\inf_abs0_m[11] ), .B(
        \un18_next_int_m[11] ), .Y(\un1_next_int[11] ));
    DFN1C0 \integ[12]  (.D(ADD_26x26_fast_I242_Y), .CLK(clk_c), .CLR(
        n_rst_c), .Q(LED_15[5]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I109_Y (.A(N427), .B(N431), .Y(
        N480));
    NOR2 \state_1_RNIVPHM[0]  (.A(\state[1]_net_1 ), .B(
        \state_1[0]_net_1 ), .Y(N_46_1));
    OA1B un1_integ_0_0_ADD_26x26_fast_I205_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\integ[22]_net_1 ), .C(\state_0[0]_net_1 ), .Y(
        ADD_26x26_fast_I205_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I115_Y (.A(N433), .B(N437), .Y(
        N486));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I12_G0N (.A(LED_15[5]), .B(
        \state[1]_net_1 ), .Y(N353));
    OR2 un1_integ_0_0_ADD_26x26_fast_I208_Y_0 (.A(N455), .B(N463), .Y(
        ADD_26x26_fast_I208_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I111_Y (.A(N433), .B(N429), .Y(
        N482));
    NOR2B \state_RNIRF7N[0]  (.A(avg_new[8]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[8] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I2_P0N (.A(\un1_next_int[2] ), .B(
        average[2]), .Y(N324));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I250_Y_0 (.A(\integ[20]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I250_Y_0));
    NOR2A \state_RNI010O[1]  (.A(\state[1]_net_1 ), .B(avg_old[8]), .Y(
        \un18_next_int_m[8] ));
    DFN1C0 \integ[10]  (.D(ADD_26x26_fast_I240_Y), .CLK(clk_c), .CLR(
        n_rst_c), .Q(LED_15[3]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I188_un1_Y (.A(N522), .B(N537), 
        .Y(I188_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I180_un1_Y (.A(N514), .B(N529), 
        .Y(I180_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I162_Y (.A(I162_un1_Y), .B(N487), 
        .Y(N541));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I6_G0N (.A(\un1_next_int[6] ), 
        .B(average[6]), .Y(N335));
    AX1D un1_integ_0_0_ADD_26x26_fast_I249_Y (.A(I180_un1_Y), .B(
        ADD_26x26_fast_I210_Y_1), .C(ADD_26x26_fast_I249_Y_0), .Y(
        \un1_integ[19] ));
    GND GND_i (.Y(GND));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I212_un1_Y_0 (.A(N480), .B(N488)
        , .C(N442), .Y(ADD_26x26_fast_I212_un1_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I1_G0N (.A(\un1_next_int[1] ), 
        .B(\integ[1]_net_1 ), .Y(N320));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I107_Y (.A(N425), .B(N429), .Y(
        N478));
    OA1B un1_integ_0_0_ADD_26x26_fast_I38_Y (.A(\integ[18]_net_1 ), .B(
        \integ[17]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N406));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I209_un1_Y_0 (.A(N512), .B(N528)
        , .Y(ADD_26x26_fast_I209_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I205_Y_3 (.A(N504), .B(N519), .C(
        ADD_26x26_fast_I205_Y_2), .Y(ADD_26x26_fast_I205_Y_3));
    AX1D un1_integ_0_0_ADD_26x26_fast_I255_Y (.A(I204_un1_Y), .B(
        ADD_26x26_fast_I204_Y_3), .C(ADD_26x26_fast_I255_Y_0), .Y(
        \un1_integ[25] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I204_Y_0 (.A(\integ[24]_net_1 ), 
        .B(\integ[23]_net_1 ), .C(\state_0[0]_net_1 ), .Y(
        ADD_26x26_fast_I204_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I243_Y (.A(N643), .B(
        ADD_26x26_fast_I243_Y_0), .Y(\un1_integ[13] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I69_Y (.A(N327), .B(N324), .Y(
        N437));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I62_Y (.A(N332), .B(average[6]), 
        .C(\un1_next_int[6] ), .Y(N430));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I193_un1_Y (.A(N478), .B(N486), 
        .C(N493), .Y(I193_un1_Y));
    NOR2A \state_RNIRRVN[1]  (.A(\state[1]_net_1 ), .B(avg_old[3]), .Y(
        \un18_next_int_m[3] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I152_un1_Y (.A(N483), .B(N476), 
        .Y(I152_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I7_G0N (.A(\un1_next_int[7] ), 
        .B(LED_15[0]), .Y(N338));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I49_Y (.A(N357), .B(N354), .Y(
        N417));
    AO1A un1_integ_0_0_ADD_26x26_fast_I42_Y (.A(\state_1[0]_net_1 ), 
        .B(\integ[16]_net_1 ), .C(N362), .Y(N410));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I145_Y (.A(N468), .B(N476), .Y(
        N522));
    OR2 un1_integ_0_0_ADD_26x26_fast_I10_P0N (.A(\un1_next_int[10] ), 
        .B(LED_15[3]), .Y(N348));
    NOR2B \state_1_RNILC4G[0]  (.A(avg_new[11]), .B(\state_1[0]_net_1 )
        , .Y(\inf_abs0_m[11] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I1_P0N (.A(\un1_next_int[1] ), .B(
        \integ[1]_net_1 ), .Y(N321));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I184_un1_Y (.A(N472), .B(N464), 
        .C(N533), .Y(I184_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I192_un1_Y (.A(N476), .B(N484), 
        .C(N491), .Y(I192_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I93_Y (.A(N363), .B(N366), .C(
        N415), .Y(N464));
    AO1B un1_integ_0_0_ADD_26x26_fast_I37_Y (.A(\integ[18]_net_1 ), .B(
        \integ[19]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N405));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I0_G0N (.A(\integ[0]_net_1 ), 
        .B(\state[1]_net_1 ), .Y(N317));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I73_Y (.A(N318), .B(N321), .Y(
        N441));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I59_Y (.A(N342), .B(N339), .Y(
        N427));
    AO1 un1_integ_0_0_ADD_26x26_fast_I52_Y (.A(N347), .B(N351), .C(
        N350), .Y(N420));
    NOR2A \state_RNO[1]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 ), 
        .Y(\state_RNO_7[1] ));
    NOR2A \state_RNI120O[1]  (.A(\state[1]_net_1 ), .B(avg_old[9]), .Y(
        \un18_next_int_m[9] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I34_Y (.A(\integ[19]_net_1 ), .B(
        \integ[20]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N402));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I236_Y (.A(\un1_next_int[6] ), 
        .B(average[6]), .C(N539), .Y(ADD_26x26_fast_I236_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I127_Y_1 (.A(
        ADD_26x26_fast_I127_Y_0), .B(N401), .Y(ADD_26x26_fast_I127_Y_1)
        );
    NOR2A \state_RNITTVN[1]  (.A(\state[1]_net_1 ), .B(avg_old[5]), .Y(
        \un18_next_int_m[5] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I150_Y (.A(I150_un1_Y), .B(N473), 
        .Y(N527));
    DFN1C0 \integ[0]  (.D(ADD_26x26_fast_I230_Y_2), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\integ[0]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I120_Y (.A(I120_un1_Y), .B(N438), 
        .Y(N491));
    AO1 un1_integ_0_0_ADD_26x26_fast_I104_Y (.A(N426), .B(N423), .C(
        N422), .Y(N475));
    NOR2A \state_RNIOOVN[1]  (.A(\state[1]_net_1 ), .B(avg_old[0]), .Y(
        \un18_next_int_m[0] ));
    VCC VCC_i (.Y(VCC));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I129_Y (.A(N399), .B(N403), .C(
        N460), .Y(N506));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I113_Y (.A(N435), .B(N431), .Y(
        N484));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I241_Y_0 (.A(\un1_next_int[11] ), 
        .B(LED_15[4]), .Y(ADD_26x26_fast_I241_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I89_Y (.A(N363), .B(N366), .C(
        N407), .Y(N460));
    AO1 un1_integ_0_0_ADD_26x26_fast_I68_Y (.A(N323), .B(N327), .C(
        N326), .Y(N436));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_0 (.A(N469), .B(N462), .C(
        N461), .Y(ADD_26x26_fast_I211_Y_0));
    NOR2A \state_RNIQQVN[1]  (.A(\state[1]_net_1 ), .B(avg_old[2]), .Y(
        \un18_next_int_m[2] ));
    DFN1C0 \integ[4]  (.D(ADD_26x26_fast_I234_Y_0_0), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(average[4]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I108_Y (.A(N430), .B(N427), .C(
        N426), .Y(N479));
    NOR2B \state_RNIQE7N[0]  (.A(avg_new[7]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[7] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I3_G0N (.A(\un18_next_int_m[3] ), 
        .B(\inf_abs0_m[3] ), .C(average[3]), .Y(N326));
    AO1 un1_integ_0_0_ADD_26x26_fast_I48_Y (.A(N353), .B(N357), .C(
        N356), .Y(N416));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I195_un1_Y (.A(N482), .B(N490), 
        .C(\un1_next_int[0] ), .Y(I195_un1_Y));
    DFN1C0 \integ[3]  (.D(ADD_26x26_fast_I233_Y_0_0), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(average[3]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I252_Y (.A(I207_un1_Y), .B(
        ADD_26x26_fast_I207_Y_2), .C(ADD_26x26_fast_I252_Y_0), .Y(
        \un1_integ[22] ));
    DFN1C0 \integ[6]  (.D(ADD_26x26_fast_I236_Y), .CLK(clk_c), .CLR(
        n_rst_c), .Q(average[6]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_1 (.A(
        ADD_26x26_fast_I210_un1_Y_0), .B(N491), .C(
        ADD_26x26_fast_I210_Y_0), .Y(ADD_26x26_fast_I210_Y_1));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y (.A(N533), .B(I194_un1_Y), 
        .C(ADD_26x26_fast_I239_Y_0), .Y(ADD_26x26_fast_I239_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I58_Y (.A(N338), .B(N342), .C(
        N341), .Y(N426));
    NOR2A \state_RNISSVN[1]  (.A(\state[1]_net_1 ), .B(avg_old[4]), .Y(
        \un18_next_int_m[4] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I67_Y (.A(average[4]), .B(
        \un1_next_int[4] ), .C(N327), .Y(N435));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I253_Y_0 (.A(\integ[23]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I253_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I64_Y (.A(N329), .B(N333), .C(
        N332), .Y(N432));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I204_un1_Y_0 (.A(N472), .B(N464)
        , .C(N502), .Y(ADD_26x26_fast_I204_un1_Y_0));
    OR2 \state_1_RNITQNB1[0]  (.A(\inf_abs0_m[10] ), .B(
        \un18_next_int_m[10] ), .Y(\un1_next_int[10] ));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I212_un1_Y (.A(N472), .B(N464), 
        .C(ADD_26x26_fast_I212_un1_Y_0), .Y(I212_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I127_Y (.A(
        ADD_26x26_fast_I127_Y_1), .B(N458), .Y(N504));
    AO1 un1_integ_0_0_ADD_26x26_fast_I110_Y (.A(N432), .B(N429), .C(
        N428), .Y(N481));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I211_un1_Y_0 (.A(N478), .B(N486)
        , .C(N493), .Y(ADD_26x26_fast_I211_un1_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I90_Y (.A(N412), .B(N408), .Y(
        N461));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I233_Y (.A(
        ADD_26x26_fast_I233_Y_0), .B(N491), .Y(
        ADD_26x26_fast_I233_Y_0_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I47_Y (.A(N360), .B(N357), .Y(
        N415));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I119_Y (.A(N441), .B(N437), .Y(
        N490));
    AO1 un1_integ_0_0_ADD_26x26_fast_I70_Y (.A(N320), .B(N324), .C(
        N323), .Y(N438));
    DFN1C0 \integ[5]  (.D(ADD_26x26_fast_I235_Y), .CLK(clk_c), .CLR(
        n_rst_c), .Q(average[5]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I182_un1_Y (.A(N516), .B(N531), 
        .Y(I182_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I161_Y (.A(N486), .B(N493), .C(
        N485), .Y(N539));
    OR2 un1_integ_0_0_ADD_26x26_fast_I44_Y (.A(N359), .B(N362), .Y(
        N412));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I245_Y (.A(N637), .B(
        ADD_26x26_fast_I245_Y_0), .Y(\un1_integ[15] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I95_Y (.A(N417), .B(N413), .Y(
        N466));
    AX1D un1_integ_0_0_ADD_26x26_fast_I239_Y_0 (.A(
        \un18_next_int_m[9] ), .B(\inf_abs0_m[9] ), .C(LED_15[2]), .Y(
        ADD_26x26_fast_I239_Y_0));
    DFN1C0 \integ[2]  (.D(ADD_26x26_fast_I232_Y_0_0), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(average[2]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I135_Y (.A(N458), .B(N466), .Y(
        N512));
    OR2 un1_integ_0_0_ADD_26x26_fast_I88_Y (.A(N410), .B(N406), .Y(
        N459));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I247_Y (.A(\state_0[0]_net_1 ), 
        .B(\integ[17]_net_1 ), .C(N633), .Y(\un1_integ[17] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I237_Y_0 (.A(LED_15[0]), .B(
        \un1_next_int[7] ), .Y(ADD_26x26_fast_I237_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I143_Y (.A(N466), .B(N474), .Y(
        N520));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I57_Y (.A(N342), .B(N345), .Y(
        N425));
    DFN1E0C0 \integ[23]  (.D(\un1_integ[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(\integ[23]_net_1 ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I8_P0N (.A(\inf_abs0_m[8] ), .B(
        \un18_next_int_m[8] ), .C(LED_15[1]), .Y(N342));
    OR3 un1_integ_0_0_ADD_26x26_fast_I212_Y (.A(I212_un1_Y), .B(N517), 
        .C(I184_un1_Y), .Y(N633));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_2 (.A(N506), .B(N521), .C(
        ADD_26x26_fast_I206_Y_1), .Y(ADD_26x26_fast_I206_Y_2));
    AO1 un1_integ_0_0_ADD_26x26_fast_I54_Y (.A(N344), .B(N348), .C(
        N347), .Y(N422));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I131_Y (.A(N401), .B(N405), .C(
        N462), .Y(N508));
    OR2A un1_integ_0_0_ADD_26x26_fast_I14_P0N (.A(\state[0]_net_1 ), 
        .B(LED_15[7]), .Y(N360));
    AX1D un1_integ_0_0_ADD_26x26_fast_I254_Y (.A(I205_un1_Y), .B(
        ADD_26x26_fast_I205_Y_3), .C(ADD_26x26_fast_I254_Y_0), .Y(
        \un1_integ[24] ));
    NOR2A un1_integ_0_0_ADD_26x26_fast_I13_G0N (.A(LED_15[6]), .B(
        \state_1[0]_net_1 ), .Y(N356));
    DFN1E0C0 \integ[19]  (.D(\un1_integ[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(\integ[19]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I117_Y (.A(N439), .B(N435), .Y(
        N488));
    DFN1E0C0 \integ[17]  (.D(\un1_integ[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(\integ[17]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I33_Y (.A(\integ[21]_net_1 ), .B(
        \integ[20]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N401));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I255_Y_0 (.A(\integ[25]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I255_Y_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I127_Y_0 (.A(\integ[22]_net_1 ), 
        .B(\integ[23]_net_1 ), .C(\state_0[0]_net_1 ), .Y(
        ADD_26x26_fast_I127_Y_0));
    DFN1E0C0 \integ[14]  (.D(\un1_integ[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(LED_15[7]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I87_Y (.A(N405), .B(N409), .Y(
        N458));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y_0 (.A(average[2]), .B(
        \un1_next_int[2] ), .Y(ADD_26x26_fast_I232_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I84_Y (.A(N406), .B(N402), .Y(
        N455));
    AO1 un1_integ_0_0_ADD_26x26_fast_I154_Y (.A(N485), .B(N478), .C(
        N477), .Y(N531));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I11_G0N (.A(\un1_next_int[11] ), 
        .B(LED_15[4]), .Y(N350));
    AO1 un1_integ_0_0_ADD_26x26_fast_I140_Y (.A(N471), .B(N464), .C(
        N463), .Y(N517));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I149_Y (.A(N472), .B(N480), .Y(
        N526));
    AO1 un1_integ_0_0_ADD_26x26_fast_I158_Y (.A(N489), .B(N482), .C(
        N481), .Y(N535));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I249_Y_0 (.A(\integ[19]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I249_Y_0));
    DFN1E0C0 \integ[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(\integ[25]_net_1 ));
    AO1 \state_0_RNIQETB1[0]  (.A(avg_new[0]), .B(\state_0[0]_net_1 ), 
        .C(\un18_next_int_m[0] ), .Y(\un1_next_int[0] ));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I242_Y (.A(\state[1]_net_1 ), .B(
        LED_15[5]), .C(N646), .Y(ADD_26x26_fast_I242_Y));
    NOR2A \state_RNIVVVN[1]  (.A(\state[1]_net_1 ), .B(avg_old[7]), .Y(
        \un18_next_int_m[7] ));
    DFN1E0C0 \integ[11]  (.D(\un1_integ[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(LED_15[4]));
    DFN1E0C0 \integ[16]  (.D(\un1_integ[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(\integ[16]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_1 (.A(
        ADD_26x26_fast_I211_un1_Y_0), .B(N516), .C(
        ADD_26x26_fast_I211_Y_0), .Y(ADD_26x26_fast_I211_Y_1));
    OR2 un1_integ_0_0_ADD_26x26_fast_I189_Y (.A(N523), .B(I189_un1_Y), 
        .Y(N640));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I254_Y_0 (.A(\integ[24]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(ADD_26x26_fast_I254_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I163_Y (.A(I163_un1_Y), .B(N489), 
        .Y(N543));
    AO1 un1_integ_0_0_ADD_26x26_fast_I96_Y (.A(N418), .B(N415), .C(
        N414), .Y(N467));
    NOR2B \state_RNINB7N[0]  (.A(avg_new[4]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[4] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I207_un1_Y (.A(
        ADD_26x26_fast_I207_un1_Y_0), .B(N539), .Y(I207_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I2_G0N (.A(\un1_next_int[2] ), 
        .B(average[2]), .Y(N323));
    AO1 un1_integ_0_0_ADD_26x26_fast_I114_Y (.A(N436), .B(N433), .C(
        N432), .Y(N485));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I189_un1_Y (.A(N478), .B(N470), 
        .C(N539), .Y(I189_un1_Y));
    DFN1C0 \integ[9]  (.D(ADD_26x26_fast_I239_Y), .CLK(clk_c), .CLR(
        n_rst_c), .Q(LED_15[2]));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I235_Y (.A(
        ADD_26x26_fast_I235_Y_0), .B(N541), .Y(ADD_26x26_fast_I235_Y));
    OA1 un1_integ_0_0_ADD_26x26_fast_I63_Y (.A(average[6]), .B(
        \un1_next_int[6] ), .C(N333), .Y(N431));
    AO1 un1_integ_0_0_ADD_26x26_fast_I118_Y (.A(N440), .B(N437), .C(
        N436), .Y(N489));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I237_Y (.A(
        ADD_26x26_fast_I237_Y_0), .B(N537), .Y(ADD_26x26_fast_I237_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I133_Y (.A(N456), .B(N464), .Y(
        N510));
    OA1B un1_integ_0_0_ADD_26x26_fast_I30_Y (.A(\integ[22]_net_1 ), .B(
        \integ[21]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N398));
    DFN1E0C0 \integ[22]  (.D(\un1_integ[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(\integ[22]_net_1 ));
    OR2 \state_RNID27F1[0]  (.A(\inf_abs0_m[1] ), .B(
        \un18_next_int_m[1] ), .Y(\un1_next_int[1] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I192_Y (.A(N529), .B(I192_un1_Y), 
        .Y(N649));
    DFN1C0 \integ[1]  (.D(ADD_26x26_fast_I231_Y_0), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\integ[1]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I35_Y (.A(\integ[20]_net_1 ), .B(
        \integ[19]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N403));
    DFN1C0 \state_0[0]  (.D(\state_1_RNIDTBQ[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_0[0]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I53_Y (.A(N351), .B(N348), .Y(
        N421));
    AO1 un1_integ_0_0_ADD_26x26_fast_I160_Y (.A(N484), .B(N491), .C(
        N483), .Y(N537));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I91_Y (.A(N409), .B(N413), .Y(
        N462));
    AX1D un1_integ_0_0_ADD_26x26_fast_I250_Y (.A(I178_un1_Y), .B(
        ADD_26x26_fast_I209_Y_1), .C(ADD_26x26_fast_I250_Y_0), .Y(
        \un1_integ[20] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I240_Y_0 (.A(LED_15[3]), .B(
        \un1_next_int[10] ), .Y(ADD_26x26_fast_I240_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I210_Y_0 (.A(N467), .B(N460), .C(
        N459), .Y(ADD_26x26_fast_I210_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I71_Y (.A(N321), .B(N324), .Y(
        N439));
    INV \integ_RNI08AC[12]  (.A(LED_15[5]), .Y(LED_15_i_0));
    DFN1E0C0 \integ[20]  (.D(\un1_integ[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(\integ[20]_net_1 ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I244_Y (.A(N640), .B(
        ADD_26x26_fast_I244_Y_0), .Y(\un1_integ[14] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I207_Y_1 (.A(N400), .B(N404), .C(
        N461), .Y(ADD_26x26_fast_I207_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I106_Y (.A(N428), .B(N425), .C(
        N424), .Y(N477));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_1 (.A(
        ADD_26x26_fast_I208_un1_Y_0), .B(N541), .C(
        ADD_26x26_fast_I208_Y_0), .Y(ADD_26x26_fast_I208_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I102_Y (.A(N424), .B(N421), .C(
        N420), .Y(N473));
    NOR2B \state_RNIOC7N[0]  (.A(avg_new[5]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[5] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I251_Y (.A(I176_un1_Y), .B(
        ADD_26x26_fast_I208_Y_1), .C(ADD_26x26_fast_I251_Y_0), .Y(
        \un1_integ[21] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I121_un1_Y (.A(N441), .B(
        \un1_next_int[0] ), .Y(I121_un1_Y));
    NOR2A un1_integ_0_0_ADD_26x26_fast_I15_G0N (.A(\integ[15]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(N362));
    DFN1E0C0 \integ[18]  (.D(\un1_integ[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(\integ[18]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I144_Y (.A(N475), .B(N468), .C(
        N467), .Y(N521));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I139_Y (.A(N462), .B(N470), .Y(
        N516));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_0 (.A(N465), .B(N458), .C(
        N457), .Y(ADD_26x26_fast_I209_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I148_Y (.A(I148_un1_Y), .B(N471), 
        .Y(N525));
    AO1 un1_integ_0_0_ADD_26x26_fast_I60_Y (.A(N335), .B(N339), .C(
        N338), .Y(N428));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y (.A(
        ADD_26x26_fast_I232_Y_0), .B(N493), .Y(
        ADD_26x26_fast_I232_Y_0_0));
    OR3 un1_integ_0_0_ADD_26x26_fast_I204_Y_2 (.A(N398), .B(
        ADD_26x26_fast_I204_Y_0), .C(N455), .Y(ADD_26x26_fast_I204_Y_2)
        );
    DFN1C0 \state[1]  (.D(\state_RNO_7[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[1]_net_1 ));
    NOR2B \state_RNIMA7N[0]  (.A(avg_new[3]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[3] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I9_G0N (.A(\un18_next_int_m[9] ), 
        .B(\inf_abs0_m[9] ), .C(LED_15[2]), .Y(N344));
    NOR2A \state_RNI9FJR[1]  (.A(\state[1]_net_1 ), .B(avg_old[10]), 
        .Y(\un18_next_int_m[10] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I40_Y (.A(\integ[17]_net_1 ), .B(
        \integ[16]_net_1 ), .C(\state_1[0]_net_1 ), .Y(N408));
    OA1 un1_integ_0_0_ADD_26x26_fast_I65_Y (.A(average[4]), .B(
        \un1_next_int[4] ), .C(N333), .Y(N433));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I207_un1_Y_0 (.A(N478), .B(N470)
        , .C(N508), .Y(ADD_26x26_fast_I207_un1_Y_0));
    NOR2B \state_RNIPD7N[0]  (.A(avg_new[6]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[6] ));
    NOR2A \state_RNIPPVN[1]  (.A(\state[1]_net_1 ), .B(avg_old[1]), .Y(
        \un18_next_int_m[1] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I188_Y (.A(N521), .B(I188_un1_Y), 
        .Y(N637));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I178_un1_Y (.A(N512), .B(N527), 
        .Y(I178_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I45_Y (.A(N360), .B(N363), .Y(
        N413));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I137_Y (.A(N460), .B(N468), .Y(
        N514));
    OR3 un1_integ_0_0_ADD_26x26_fast_I3_P0N (.A(\un18_next_int_m[3] ), 
        .B(\inf_abs0_m[3] ), .C(average[3]), .Y(N327));
    AX1D un1_integ_0_0_ADD_26x26_fast_I233_Y_0 (.A(
        \un18_next_int_m[3] ), .B(\inf_abs0_m[3] ), .C(average[3]), .Y(
        ADD_26x26_fast_I233_Y_0));
    OR2A un1_integ_0_0_ADD_26x26_fast_I16_P0N (.A(\state_1[0]_net_1 ), 
        .B(\integ[16]_net_1 ), .Y(N366));
    AO1 un1_integ_0_0_ADD_26x26_fast_I50_Y (.A(N350), .B(N354), .C(
        N353), .Y(N418));
    AO1 un1_integ_0_0_ADD_26x26_fast_I204_Y_3 (.A(N502), .B(N517), .C(
        ADD_26x26_fast_I204_Y_2), .Y(ADD_26x26_fast_I204_Y_3));
    OR2 \state_RNINC7F1[0]  (.A(\inf_abs0_m[6] ), .B(
        \un18_next_int_m[6] ), .Y(\un1_next_int[6] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I36_Y (.A(\integ[18]_net_1 ), .B(
        \integ[19]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N404));
    NOR2A \state_RNIUUVN[1]  (.A(\state[1]_net_1 ), .B(avg_old[6]), .Y(
        \un18_next_int_m[6] ));
    NOR2B \state_RNISG7N[0]  (.A(avg_new[9]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[9] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I0_P0N (.A(\integ[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(N318));
    OR2 \state_RNIF47F1[0]  (.A(\inf_abs0_m[2] ), .B(
        \un18_next_int_m[2] ), .Y(\un1_next_int[2] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I55_Y (.A(N348), .B(N345), .Y(
        N423));
    NOR2B \state_1_RNIDTBQ[0]  (.A(N_46_1), .B(calc_avg), .Y(
        \state_1_RNIDTBQ[0]_net_1 ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I205_un1_Y (.A(N535), .B(
        I195_un1_Y), .C(ADD_26x26_fast_I205_un1_Y_0), .Y(I205_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I163_un1_Y (.A(N490), .B(
        \un1_next_int[0] ), .Y(I163_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I120_un1_Y (.A(N439), .B(N442), 
        .Y(I120_un1_Y));
    OR3 un1_integ_0_0_ADD_26x26_fast_I206_Y_1 (.A(N402), .B(N398), .C(
        N459), .Y(ADD_26x26_fast_I206_Y_1));
    OA1 un1_integ_0_0_ADD_26x26_fast_I5_G0N (.A(\un18_next_int_m[5] ), 
        .B(\inf_abs0_m[5] ), .C(average[5]), .Y(N332));
    DFN1C0 \integ[7]  (.D(ADD_26x26_fast_I237_Y), .CLK(clk_c), .CLR(
        n_rst_c), .Q(LED_15[0]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_2 (.A(N508), .B(N523), .C(
        ADD_26x26_fast_I207_Y_1), .Y(ADD_26x26_fast_I207_Y_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I4_G0N (.A(\un1_next_int[4] ), 
        .B(average[4]), .Y(N329));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y (.A(
        ADD_26x26_fast_I234_Y_0), .B(N543), .Y(
        ADD_26x26_fast_I234_Y_0_0));
    OR3 un1_integ_0_0_ADD_26x26_fast_I205_Y_2 (.A(N400), .B(
        ADD_26x26_fast_I205_Y_0), .C(N457), .Y(ADD_26x26_fast_I205_Y_2)
        );
    NOR2B un1_integ_0_0_ADD_26x26_fast_I162_un1_Y (.A(N488), .B(N442), 
        .Y(I162_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I240_Y (.A(N531), .B(I193_un1_Y), 
        .C(ADD_26x26_fast_I240_Y_0), .Y(ADD_26x26_fast_I240_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I156_Y (.A(N487), .B(N480), .C(
        N479), .Y(N533));
    DFN1C0 \integ[8]  (.D(ADD_26x26_fast_I238_Y), .CLK(clk_c), .CLR(
        n_rst_c), .Q(LED_15[1]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I85_Y (.A(N403), .B(N407), .Y(
        N456));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I251_Y_0 (.A(\integ[21]_net_1 ), 
        .B(\state_1[0]_net_1 ), .Y(ADD_26x26_fast_I251_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I152_Y (.A(I152_un1_Y), .B(N475), 
        .Y(N529));
    OR3 un1_integ_0_0_ADD_26x26_fast_I9_P0N (.A(\un18_next_int_m[9] ), 
        .B(\inf_abs0_m[9] ), .C(LED_15[2]), .Y(N345));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I208_un1_Y_0 (.A(N510), .B(N526)
        , .Y(ADD_26x26_fast_I208_un1_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I191_Y (.A(N528), .B(N543), .C(
        N527), .Y(N646));
    AO1B un1_integ_0_0_ADD_26x26_fast_I31_Y (.A(\integ[22]_net_1 ), .B(
        \integ[21]_net_1 ), .C(\state_0[0]_net_1 ), .Y(N399));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I206_un1_Y (.A(N522), .B(N506), 
        .C(N537), .Y(I206_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I235_Y_0 (.A(
        \un18_next_int_m[5] ), .B(\inf_abs0_m[5] ), .C(average[5]), .Y(
        ADD_26x26_fast_I235_Y_0));
    NOR2B \state_1_RNIKB4G[0]  (.A(avg_new[10]), .B(\state_1[0]_net_1 )
        , .Y(\inf_abs0_m[10] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I241_Y (.A(N649), .B(
        ADD_26x26_fast_I241_Y_0), .Y(\un1_integ[11] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I11_P0N (.A(\un1_next_int[11] ), 
        .B(LED_15[4]), .Y(N351));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I243_Y_0 (.A(LED_15[6]), .B(
        \state[0]_net_1 ), .Y(ADD_26x26_fast_I243_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I105_Y (.A(N423), .B(N427), .Y(
        N476));
    AO1 un1_integ_0_0_ADD_26x26_fast_I213_Y_0 (.A(
        ADD_26x26_fast_I213_un1_Y_0), .B(N520), .C(N519), .Y(
        ADD_26x26_fast_I213_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I238_Y_0 (.A(\inf_abs0_m[8] ), 
        .B(\un18_next_int_m[8] ), .C(LED_15[1]), .Y(
        ADD_26x26_fast_I238_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I101_Y (.A(N423), .B(N419), .Y(
        N472));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I66_Y (.A(N326), .B(average[4]), 
        .C(\un1_next_int[4] ), .Y(N434));
    AX1D un1_integ_0_0_ADD_26x26_fast_I248_Y (.A(I182_un1_Y), .B(
        ADD_26x26_fast_I211_Y_1), .C(ADD_26x26_fast_I248_Y_0), .Y(
        \un1_integ[18] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I99_Y (.A(N417), .B(N421), .Y(
        N470));
    OR2 un1_integ_0_0_ADD_26x26_fast_I92_Y (.A(N414), .B(N410), .Y(
        N463));
    AO1 un1_integ_0_0_ADD_26x26_fast_I72_Y (.A(N317), .B(N321), .C(
        N320), .Y(N440));
    OR2A un1_integ_0_0_ADD_26x26_fast_I13_P0N (.A(\state_1[0]_net_1 ), 
        .B(LED_15[6]), .Y(N357));
    OR2 un1_integ_0_0_ADD_26x26_fast_I46_Y (.A(N356), .B(N359), .Y(
        N414));
    NOR2B \state_RNIL97N[0]  (.A(avg_new[2]), .B(\state[0]_net_1 ), .Y(
        \inf_abs0_m[2] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I116_Y (.A(N438), .B(N435), .C(
        N434), .Y(N487));
    AO1 un1_integ_0_0_ADD_26x26_fast_I112_Y (.A(N434), .B(N431), .C(
        N430), .Y(N483));
    OR2 \state_RNIPE7F1[0]  (.A(\inf_abs0_m[7] ), .B(
        \un18_next_int_m[7] ), .Y(\un1_next_int[7] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I8_G0N (.A(\inf_abs0_m[8] ), .B(
        \un18_next_int_m[8] ), .C(LED_15[1]), .Y(N341));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I213_un1_Y_0 (.A(N482), .B(N490)
        , .C(\un1_next_int[0] ), .Y(ADD_26x26_fast_I213_un1_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y_0 (.A(average[4]), .B(
        \un1_next_int[4] ), .Y(ADD_26x26_fast_I234_Y_0));
    
endmodule


module error_sr_13s_5s_3(
       cur_vd,
       avg_new,
       avg_old,
       avg_enable_0,
       avg_enable,
       avg_enable_1,
       n_rst_c,
       clk_c
    );
input  [11:0] cur_vd;
output [11:0] avg_new;
output [11:0] avg_old;
input  avg_enable_0;
input  avg_enable;
input  avg_enable_1;
input  n_rst_c;
input  clk_c;

    wire \sr_3_[0]_net_1 , \sr_3_[1]_net_1 , \sr_3_[2]_net_1 , 
        \sr_3_[3]_net_1 , \sr_3_[4]_net_1 , \sr_3_[5]_net_1 , 
        \sr_3_[6]_net_1 , \sr_3_[7]_net_1 , \sr_3_[8]_net_1 , 
        \sr_3_[9]_net_1 , \sr_3_[10]_net_1 , \sr_3_[11]_net_1 , 
        \sr_2_[0]_net_1 , \sr_2_[1]_net_1 , \sr_2_[2]_net_1 , 
        \sr_2_[3]_net_1 , \sr_2_[4]_net_1 , \sr_2_[5]_net_1 , 
        \sr_2_[6]_net_1 , \sr_2_[7]_net_1 , \sr_2_[8]_net_1 , 
        \sr_2_[9]_net_1 , \sr_2_[10]_net_1 , \sr_2_[11]_net_1 , 
        \sr_1_[0]_net_1 , \sr_1_[1]_net_1 , \sr_1_[2]_net_1 , 
        \sr_1_[3]_net_1 , \sr_1_[4]_net_1 , \sr_1_[5]_net_1 , 
        \sr_1_[6]_net_1 , \sr_1_[7]_net_1 , \sr_1_[8]_net_1 , 
        \sr_1_[9]_net_1 , \sr_1_[10]_net_1 , \sr_1_[11]_net_1 , GND, 
        VCC;
    
    DFN1E1C0 \sr_1_[11]  (.D(avg_new[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[11]_net_1 ));
    DFN1E1C0 \sr_3_[3]  (.D(\sr_2_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_3_[3]_net_1 ));
    DFN1E1C0 \sr_4_[4]  (.D(\sr_3_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[4]));
    DFN1E1C0 \sr_0_[10]  (.D(cur_vd[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(avg_new[10]));
    DFN1E1C0 \sr_4_[8]  (.D(\sr_3_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[8]));
    DFN1E1C0 \sr_4_[0]  (.D(\sr_3_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(avg_old[0]));
    DFN1E1C0 \sr_1_[2]  (.D(avg_new[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable), .Q(\sr_1_[2]_net_1 ));
    DFN1E1C0 \sr_0_[2]  (.D(cur_vd[2]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[2]));
    DFN1E1C0 \sr_2_[2]  (.D(\sr_1_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[2]_net_1 ));
    DFN1E1C0 \sr_0_[11]  (.D(cur_vd[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(avg_new[11]));
    DFN1E1C0 \sr_1_[3]  (.D(avg_new[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable), .Q(\sr_1_[3]_net_1 ));
    DFN1E1C0 \sr_0_[3]  (.D(cur_vd[3]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[3]));
    DFN1E1C0 \sr_1_[10]  (.D(avg_new[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable_0), .Q(\sr_1_[10]_net_1 ));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \sr_4_[10]  (.D(\sr_3_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[10]));
    DFN1E1C0 \sr_3_[11]  (.D(\sr_2_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_3_[11]_net_1 ));
    DFN1E1C0 \sr_2_[3]  (.D(\sr_1_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[3]_net_1 ));
    DFN1E1C0 \sr_3_[6]  (.D(\sr_2_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[6]_net_1 ));
    DFN1E1C0 \sr_3_[1]  (.D(\sr_2_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_3_[1]_net_1 ));
    DFN1E1C0 \sr_4_[2]  (.D(\sr_3_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(avg_old[2]));
    DFN1E1C0 \sr_1_[6]  (.D(avg_new[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable), .Q(\sr_1_[6]_net_1 ));
    DFN1E1C0 \sr_4_[3]  (.D(\sr_3_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(avg_old[3]));
    DFN1E1C0 \sr_0_[6]  (.D(cur_vd[6]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[6]));
    DFN1E1C0 \sr_3_[9]  (.D(\sr_2_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[9]_net_1 ));
    DFN1E1C0 \sr_1_[1]  (.D(avg_new[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable), .Q(\sr_1_[1]_net_1 ));
    DFN1E1C0 \sr_0_[1]  (.D(cur_vd[1]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[1]));
    DFN1E1C0 \sr_2_[6]  (.D(\sr_1_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[6]_net_1 ));
    DFN1E1C0 \sr_2_[1]  (.D(\sr_1_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[1]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1C0 \sr_3_[5]  (.D(\sr_2_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[5]_net_1 ));
    DFN1E1C0 \sr_3_[7]  (.D(\sr_2_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[7]_net_1 ));
    DFN1E1C0 \sr_1_[9]  (.D(avg_new[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable), .Q(\sr_1_[9]_net_1 ));
    DFN1E1C0 \sr_0_[9]  (.D(cur_vd[9]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[9]));
    DFN1E1C0 \sr_2_[11]  (.D(\sr_1_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[11]_net_1 ));
    DFN1E1C0 \sr_4_[6]  (.D(\sr_3_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[6]));
    DFN1E1C0 \sr_2_[9]  (.D(\sr_1_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[9]_net_1 ));
    DFN1E1C0 \sr_4_[11]  (.D(\sr_3_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[11]));
    DFN1E1C0 \sr_4_[1]  (.D(\sr_3_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(avg_old[1]));
    DFN1E1C0 \sr_3_[4]  (.D(\sr_2_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_3_[4]_net_1 ));
    DFN1E1C0 \sr_1_[5]  (.D(avg_new[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable), .Q(\sr_1_[5]_net_1 ));
    DFN1E1C0 \sr_0_[5]  (.D(cur_vd[5]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[5]));
    DFN1E1C0 \sr_1_[7]  (.D(avg_new[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable), .Q(\sr_1_[7]_net_1 ));
    DFN1E1C0 \sr_0_[7]  (.D(cur_vd[7]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[7]));
    DFN1E1C0 \sr_3_[8]  (.D(\sr_2_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_3_[8]_net_1 ));
    DFN1E1C0 \sr_3_[0]  (.D(\sr_2_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_3_[0]_net_1 ));
    DFN1E1C0 \sr_2_[5]  (.D(\sr_1_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[5]_net_1 ));
    DFN1E1C0 \sr_2_[7]  (.D(\sr_1_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[7]_net_1 ));
    DFN1E1C0 \sr_4_[9]  (.D(\sr_3_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[9]));
    DFN1E1C0 \sr_1_[4]  (.D(avg_new[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable), .Q(\sr_1_[4]_net_1 ));
    DFN1E1C0 \sr_0_[4]  (.D(cur_vd[4]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[4]));
    DFN1E1C0 \sr_1_[8]  (.D(avg_new[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable), .Q(\sr_1_[8]_net_1 ));
    DFN1E1C0 \sr_1_[0]  (.D(avg_new[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(avg_enable), .Q(\sr_1_[0]_net_1 ));
    DFN1E1C0 \sr_2_[4]  (.D(\sr_1_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[4]_net_1 ));
    DFN1E1C0 \sr_0_[8]  (.D(cur_vd[8]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[8]));
    DFN1E1C0 \sr_0_[0]  (.D(cur_vd[0]), .CLK(clk_c), .CLR(n_rst_c), .E(
        avg_enable_1), .Q(avg_new[0]));
    DFN1E1C0 \sr_4_[5]  (.D(\sr_3_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[5]));
    DFN1E1C0 \sr_2_[8]  (.D(\sr_1_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[8]_net_1 ));
    DFN1E1C0 \sr_2_[0]  (.D(\sr_1_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_2_[0]_net_1 ));
    DFN1E1C0 \sr_4_[7]  (.D(\sr_3_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable), .Q(avg_old[7]));
    DFN1E1C0 \sr_3_[10]  (.D(\sr_2_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_3_[10]_net_1 ));
    DFN1E1C0 \sr_3_[2]  (.D(\sr_2_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_0), .Q(\sr_3_[2]_net_1 ));
    DFN1E1C0 \sr_2_[10]  (.D(\sr_1_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(avg_enable_1), .Q(\sr_2_[10]_net_1 ));
    
endmodule


module error_sr_13s_64s_3(
       sr_old,
       sr_new,
       cur_error,
       sr_prev,
       sr_new_0_0,
       int_enable,
       n_rst_c,
       clk_c
    );
output [12:0] sr_old;
output [12:0] sr_new;
input  [12:0] cur_error;
output [12:0] sr_prev;
output sr_new_0_0;
input  int_enable;
input  n_rst_c;
input  clk_c;

    wire \sr_9_[0]_net_1 , \sr_8_[0]_net_1 , \sr_9_[1]_net_1 , 
        \sr_8_[1]_net_1 , \sr_9_[2]_net_1 , \sr_8_[2]_net_1 , 
        \sr_9_[3]_net_1 , \sr_8_[3]_net_1 , \sr_9_[4]_net_1 , 
        \sr_8_[4]_net_1 , \sr_9_[5]_net_1 , \sr_8_[5]_net_1 , 
        \sr_9_[6]_net_1 , \sr_8_[6]_net_1 , \sr_9_[7]_net_1 , 
        \sr_8_[7]_net_1 , \sr_9_[8]_net_1 , \sr_8_[8]_net_1 , 
        \sr_9_[9]_net_1 , \sr_8_[9]_net_1 , \sr_9_[10]_net_1 , 
        \sr_8_[10]_net_1 , \sr_9_[11]_net_1 , \sr_8_[11]_net_1 , 
        \sr_9_[12]_net_1 , \sr_8_[12]_net_1 , \sr_7_[0]_net_1 , 
        \sr_7_[1]_net_1 , \sr_7_[2]_net_1 , \sr_7_[3]_net_1 , 
        \sr_7_[4]_net_1 , \sr_7_[5]_net_1 , \sr_7_[6]_net_1 , 
        \sr_7_[7]_net_1 , \sr_7_[8]_net_1 , \sr_7_[9]_net_1 , 
        \sr_7_[10]_net_1 , \sr_7_[11]_net_1 , \sr_7_[12]_net_1 , 
        \sr_6_[0]_net_1 , \sr_6_[1]_net_1 , \sr_6_[2]_net_1 , 
        \sr_6_[3]_net_1 , \sr_6_[4]_net_1 , \sr_6_[5]_net_1 , 
        \sr_6_[6]_net_1 , \sr_6_[7]_net_1 , \sr_6_[8]_net_1 , 
        \sr_6_[9]_net_1 , \sr_6_[10]_net_1 , \sr_6_[11]_net_1 , 
        \sr_6_[12]_net_1 , \sr_5_[0]_net_1 , \sr_5_[1]_net_1 , 
        \sr_5_[2]_net_1 , \sr_5_[3]_net_1 , \sr_5_[4]_net_1 , 
        \sr_5_[5]_net_1 , \sr_5_[6]_net_1 , \sr_5_[7]_net_1 , 
        \sr_5_[8]_net_1 , \sr_5_[9]_net_1 , \sr_5_[10]_net_1 , 
        \sr_5_[11]_net_1 , \sr_5_[12]_net_1 , \sr_4_[0]_net_1 , 
        \sr_4_[1]_net_1 , \sr_4_[2]_net_1 , \sr_4_[3]_net_1 , 
        \sr_4_[4]_net_1 , \sr_4_[5]_net_1 , \sr_4_[6]_net_1 , 
        \sr_4_[7]_net_1 , \sr_4_[8]_net_1 , \sr_4_[9]_net_1 , 
        \sr_4_[10]_net_1 , \sr_4_[11]_net_1 , \sr_4_[12]_net_1 , 
        \sr_3_[0]_net_1 , \sr_3_[1]_net_1 , \sr_3_[2]_net_1 , 
        \sr_3_[3]_net_1 , \sr_3_[4]_net_1 , \sr_3_[5]_net_1 , 
        \sr_3_[6]_net_1 , \sr_3_[7]_net_1 , \sr_3_[8]_net_1 , 
        \sr_3_[9]_net_1 , \sr_3_[10]_net_1 , \sr_3_[11]_net_1 , 
        \sr_3_[12]_net_1 , \sr_2_[0]_net_1 , \sr_2_[1]_net_1 , 
        \sr_2_[2]_net_1 , \sr_2_[3]_net_1 , \sr_2_[4]_net_1 , 
        \sr_2_[5]_net_1 , \sr_2_[6]_net_1 , \sr_2_[7]_net_1 , 
        \sr_2_[8]_net_1 , \sr_2_[9]_net_1 , \sr_2_[10]_net_1 , 
        \sr_2_[11]_net_1 , \sr_2_[12]_net_1 , \sr_24_[0]_net_1 , 
        \sr_23_[0]_net_1 , \sr_24_[1]_net_1 , \sr_23_[1]_net_1 , 
        \sr_24_[2]_net_1 , \sr_23_[2]_net_1 , \sr_24_[3]_net_1 , 
        \sr_23_[3]_net_1 , \sr_24_[4]_net_1 , \sr_23_[4]_net_1 , 
        \sr_24_[5]_net_1 , \sr_23_[5]_net_1 , \sr_24_[6]_net_1 , 
        \sr_23_[6]_net_1 , \sr_24_[7]_net_1 , \sr_23_[7]_net_1 , 
        \sr_24_[8]_net_1 , \sr_23_[8]_net_1 , \sr_24_[9]_net_1 , 
        \sr_23_[9]_net_1 , \sr_24_[10]_net_1 , \sr_23_[10]_net_1 , 
        \sr_24_[11]_net_1 , \sr_23_[11]_net_1 , \sr_24_[12]_net_1 , 
        \sr_23_[12]_net_1 , \sr_22_[0]_net_1 , \sr_22_[1]_net_1 , 
        \sr_22_[2]_net_1 , \sr_22_[3]_net_1 , \sr_22_[4]_net_1 , 
        \sr_22_[5]_net_1 , \sr_22_[6]_net_1 , \sr_22_[7]_net_1 , 
        \sr_22_[8]_net_1 , \sr_22_[9]_net_1 , \sr_22_[10]_net_1 , 
        \sr_22_[11]_net_1 , \sr_22_[12]_net_1 , \sr_21_[0]_net_1 , 
        \sr_21_[1]_net_1 , \sr_21_[2]_net_1 , \sr_21_[3]_net_1 , 
        \sr_21_[4]_net_1 , \sr_21_[5]_net_1 , \sr_21_[6]_net_1 , 
        \sr_21_[7]_net_1 , \sr_21_[8]_net_1 , \sr_21_[9]_net_1 , 
        \sr_21_[10]_net_1 , \sr_21_[11]_net_1 , \sr_21_[12]_net_1 , 
        \sr_20_[0]_net_1 , \sr_20_[1]_net_1 , \sr_20_[2]_net_1 , 
        \sr_20_[3]_net_1 , \sr_20_[4]_net_1 , \sr_20_[5]_net_1 , 
        \sr_20_[6]_net_1 , \sr_20_[7]_net_1 , \sr_20_[8]_net_1 , 
        \sr_20_[9]_net_1 , \sr_20_[10]_net_1 , \sr_20_[11]_net_1 , 
        \sr_20_[12]_net_1 , \sr_19_[0]_net_1 , \sr_19_[1]_net_1 , 
        \sr_19_[2]_net_1 , \sr_19_[3]_net_1 , \sr_19_[4]_net_1 , 
        \sr_19_[5]_net_1 , \sr_19_[6]_net_1 , \sr_19_[7]_net_1 , 
        \sr_19_[8]_net_1 , \sr_19_[9]_net_1 , \sr_19_[10]_net_1 , 
        \sr_19_[11]_net_1 , \sr_19_[12]_net_1 , \sr_18_[0]_net_1 , 
        \sr_18_[1]_net_1 , \sr_18_[2]_net_1 , \sr_18_[3]_net_1 , 
        \sr_18_[4]_net_1 , \sr_18_[5]_net_1 , \sr_18_[6]_net_1 , 
        \sr_18_[7]_net_1 , \sr_18_[8]_net_1 , \sr_18_[9]_net_1 , 
        \sr_18_[10]_net_1 , \sr_18_[11]_net_1 , \sr_18_[12]_net_1 , 
        \sr_17_[0]_net_1 , \sr_17_[1]_net_1 , \sr_17_[2]_net_1 , 
        \sr_17_[3]_net_1 , \sr_17_[4]_net_1 , \sr_17_[5]_net_1 , 
        \sr_17_[6]_net_1 , \sr_17_[7]_net_1 , \sr_17_[8]_net_1 , 
        \sr_17_[9]_net_1 , \sr_17_[10]_net_1 , \sr_17_[11]_net_1 , 
        \sr_17_[12]_net_1 , \sr_16_[0]_net_1 , \sr_16_[1]_net_1 , 
        \sr_16_[2]_net_1 , \sr_16_[3]_net_1 , \sr_16_[4]_net_1 , 
        \sr_16_[5]_net_1 , \sr_16_[6]_net_1 , \sr_16_[7]_net_1 , 
        \sr_16_[8]_net_1 , \sr_16_[9]_net_1 , \sr_16_[10]_net_1 , 
        \sr_16_[11]_net_1 , \sr_16_[12]_net_1 , \sr_15_[0]_net_1 , 
        \sr_15_[1]_net_1 , \sr_15_[2]_net_1 , \sr_15_[3]_net_1 , 
        \sr_15_[4]_net_1 , \sr_15_[5]_net_1 , \sr_15_[6]_net_1 , 
        \sr_15_[7]_net_1 , \sr_15_[8]_net_1 , \sr_15_[9]_net_1 , 
        \sr_15_[10]_net_1 , \sr_15_[11]_net_1 , \sr_15_[12]_net_1 , 
        \sr_14_[0]_net_1 , \sr_14_[1]_net_1 , \sr_14_[2]_net_1 , 
        \sr_14_[3]_net_1 , \sr_14_[4]_net_1 , \sr_14_[5]_net_1 , 
        \sr_14_[6]_net_1 , \sr_14_[7]_net_1 , \sr_14_[8]_net_1 , 
        \sr_14_[9]_net_1 , \sr_14_[10]_net_1 , \sr_14_[11]_net_1 , 
        \sr_14_[12]_net_1 , \sr_13_[0]_net_1 , \sr_13_[1]_net_1 , 
        \sr_13_[2]_net_1 , \sr_13_[3]_net_1 , \sr_13_[4]_net_1 , 
        \sr_13_[5]_net_1 , \sr_13_[6]_net_1 , \sr_13_[7]_net_1 , 
        \sr_13_[8]_net_1 , \sr_13_[9]_net_1 , \sr_13_[10]_net_1 , 
        \sr_13_[11]_net_1 , \sr_13_[12]_net_1 , \sr_12_[0]_net_1 , 
        \sr_12_[1]_net_1 , \sr_12_[2]_net_1 , \sr_12_[3]_net_1 , 
        \sr_12_[4]_net_1 , \sr_12_[5]_net_1 , \sr_12_[6]_net_1 , 
        \sr_12_[7]_net_1 , \sr_12_[8]_net_1 , \sr_12_[9]_net_1 , 
        \sr_12_[10]_net_1 , \sr_12_[11]_net_1 , \sr_12_[12]_net_1 , 
        \sr_11_[0]_net_1 , \sr_11_[1]_net_1 , \sr_11_[2]_net_1 , 
        \sr_11_[3]_net_1 , \sr_11_[4]_net_1 , \sr_11_[5]_net_1 , 
        \sr_11_[6]_net_1 , \sr_11_[7]_net_1 , \sr_11_[8]_net_1 , 
        \sr_11_[9]_net_1 , \sr_11_[10]_net_1 , \sr_11_[11]_net_1 , 
        \sr_11_[12]_net_1 , \sr_10_[0]_net_1 , \sr_10_[1]_net_1 , 
        \sr_10_[2]_net_1 , \sr_10_[3]_net_1 , \sr_10_[4]_net_1 , 
        \sr_10_[5]_net_1 , \sr_10_[6]_net_1 , \sr_10_[7]_net_1 , 
        \sr_10_[8]_net_1 , \sr_10_[9]_net_1 , \sr_10_[10]_net_1 , 
        \sr_10_[11]_net_1 , \sr_10_[12]_net_1 , \sr_39_[0]_net_1 , 
        \sr_38_[0]_net_1 , \sr_39_[1]_net_1 , \sr_38_[1]_net_1 , 
        \sr_39_[2]_net_1 , \sr_38_[2]_net_1 , \sr_39_[3]_net_1 , 
        \sr_38_[3]_net_1 , \sr_39_[4]_net_1 , \sr_38_[4]_net_1 , 
        \sr_39_[5]_net_1 , \sr_38_[5]_net_1 , \sr_39_[6]_net_1 , 
        \sr_38_[6]_net_1 , \sr_39_[7]_net_1 , \sr_38_[7]_net_1 , 
        \sr_39_[8]_net_1 , \sr_38_[8]_net_1 , \sr_39_[9]_net_1 , 
        \sr_38_[9]_net_1 , \sr_39_[10]_net_1 , \sr_38_[10]_net_1 , 
        \sr_39_[11]_net_1 , \sr_38_[11]_net_1 , \sr_39_[12]_net_1 , 
        \sr_38_[12]_net_1 , \sr_37_[0]_net_1 , \sr_37_[1]_net_1 , 
        \sr_37_[2]_net_1 , \sr_37_[3]_net_1 , \sr_37_[4]_net_1 , 
        \sr_37_[5]_net_1 , \sr_37_[6]_net_1 , \sr_37_[7]_net_1 , 
        \sr_37_[8]_net_1 , \sr_37_[9]_net_1 , \sr_37_[10]_net_1 , 
        \sr_37_[11]_net_1 , \sr_37_[12]_net_1 , \sr_36_[0]_net_1 , 
        \sr_36_[1]_net_1 , \sr_36_[2]_net_1 , \sr_36_[3]_net_1 , 
        \sr_36_[4]_net_1 , \sr_36_[5]_net_1 , \sr_36_[6]_net_1 , 
        \sr_36_[7]_net_1 , \sr_36_[8]_net_1 , \sr_36_[9]_net_1 , 
        \sr_36_[10]_net_1 , \sr_36_[11]_net_1 , \sr_36_[12]_net_1 , 
        \sr_35_[0]_net_1 , \sr_35_[1]_net_1 , \sr_35_[2]_net_1 , 
        \sr_35_[3]_net_1 , \sr_35_[4]_net_1 , \sr_35_[5]_net_1 , 
        \sr_35_[6]_net_1 , \sr_35_[7]_net_1 , \sr_35_[8]_net_1 , 
        \sr_35_[9]_net_1 , \sr_35_[10]_net_1 , \sr_35_[11]_net_1 , 
        \sr_35_[12]_net_1 , \sr_34_[0]_net_1 , \sr_34_[1]_net_1 , 
        \sr_34_[2]_net_1 , \sr_34_[3]_net_1 , \sr_34_[4]_net_1 , 
        \sr_34_[5]_net_1 , \sr_34_[6]_net_1 , \sr_34_[7]_net_1 , 
        \sr_34_[8]_net_1 , \sr_34_[9]_net_1 , \sr_34_[10]_net_1 , 
        \sr_34_[11]_net_1 , \sr_34_[12]_net_1 , \sr_33_[0]_net_1 , 
        \sr_33_[1]_net_1 , \sr_33_[2]_net_1 , \sr_33_[3]_net_1 , 
        \sr_33_[4]_net_1 , \sr_33_[5]_net_1 , \sr_33_[6]_net_1 , 
        \sr_33_[7]_net_1 , \sr_33_[8]_net_1 , \sr_33_[9]_net_1 , 
        \sr_33_[10]_net_1 , \sr_33_[11]_net_1 , \sr_33_[12]_net_1 , 
        \sr_32_[0]_net_1 , \sr_32_[1]_net_1 , \sr_32_[2]_net_1 , 
        \sr_32_[3]_net_1 , \sr_32_[4]_net_1 , \sr_32_[5]_net_1 , 
        \sr_32_[6]_net_1 , \sr_32_[7]_net_1 , \sr_32_[8]_net_1 , 
        \sr_32_[9]_net_1 , \sr_32_[10]_net_1 , \sr_32_[11]_net_1 , 
        \sr_32_[12]_net_1 , \sr_31_[0]_net_1 , \sr_31_[1]_net_1 , 
        \sr_31_[2]_net_1 , \sr_31_[3]_net_1 , \sr_31_[4]_net_1 , 
        \sr_31_[5]_net_1 , \sr_31_[6]_net_1 , \sr_31_[7]_net_1 , 
        \sr_31_[8]_net_1 , \sr_31_[9]_net_1 , \sr_31_[10]_net_1 , 
        \sr_31_[11]_net_1 , \sr_31_[12]_net_1 , \sr_30_[0]_net_1 , 
        \sr_30_[1]_net_1 , \sr_30_[2]_net_1 , \sr_30_[3]_net_1 , 
        \sr_30_[4]_net_1 , \sr_30_[5]_net_1 , \sr_30_[6]_net_1 , 
        \sr_30_[7]_net_1 , \sr_30_[8]_net_1 , \sr_30_[9]_net_1 , 
        \sr_30_[10]_net_1 , \sr_30_[11]_net_1 , \sr_30_[12]_net_1 , 
        \sr_29_[0]_net_1 , \sr_29_[1]_net_1 , \sr_29_[2]_net_1 , 
        \sr_29_[3]_net_1 , \sr_29_[4]_net_1 , \sr_29_[5]_net_1 , 
        \sr_29_[6]_net_1 , \sr_29_[7]_net_1 , \sr_29_[8]_net_1 , 
        \sr_29_[9]_net_1 , \sr_29_[10]_net_1 , \sr_29_[11]_net_1 , 
        \sr_29_[12]_net_1 , \sr_28_[0]_net_1 , \sr_28_[1]_net_1 , 
        \sr_28_[2]_net_1 , \sr_28_[3]_net_1 , \sr_28_[4]_net_1 , 
        \sr_28_[5]_net_1 , \sr_28_[6]_net_1 , \sr_28_[7]_net_1 , 
        \sr_28_[8]_net_1 , \sr_28_[9]_net_1 , \sr_28_[10]_net_1 , 
        \sr_28_[11]_net_1 , \sr_28_[12]_net_1 , \sr_27_[0]_net_1 , 
        \sr_27_[1]_net_1 , \sr_27_[2]_net_1 , \sr_27_[3]_net_1 , 
        \sr_27_[4]_net_1 , \sr_27_[5]_net_1 , \sr_27_[6]_net_1 , 
        \sr_27_[7]_net_1 , \sr_27_[8]_net_1 , \sr_27_[9]_net_1 , 
        \sr_27_[10]_net_1 , \sr_27_[11]_net_1 , \sr_27_[12]_net_1 , 
        \sr_26_[0]_net_1 , \sr_26_[1]_net_1 , \sr_26_[2]_net_1 , 
        \sr_26_[3]_net_1 , \sr_26_[4]_net_1 , \sr_26_[5]_net_1 , 
        \sr_26_[6]_net_1 , \sr_26_[7]_net_1 , \sr_26_[8]_net_1 , 
        \sr_26_[9]_net_1 , \sr_26_[10]_net_1 , \sr_26_[11]_net_1 , 
        \sr_26_[12]_net_1 , \sr_25_[0]_net_1 , \sr_25_[1]_net_1 , 
        \sr_25_[2]_net_1 , \sr_25_[3]_net_1 , \sr_25_[4]_net_1 , 
        \sr_25_[5]_net_1 , \sr_25_[6]_net_1 , \sr_25_[7]_net_1 , 
        \sr_25_[8]_net_1 , \sr_25_[9]_net_1 , \sr_25_[10]_net_1 , 
        \sr_25_[11]_net_1 , \sr_25_[12]_net_1 , \sr_54_[0]_net_1 , 
        \sr_53_[0]_net_1 , \sr_54_[1]_net_1 , \sr_53_[1]_net_1 , 
        \sr_54_[2]_net_1 , \sr_53_[2]_net_1 , \sr_54_[3]_net_1 , 
        \sr_53_[3]_net_1 , \sr_54_[4]_net_1 , \sr_53_[4]_net_1 , 
        \sr_54_[5]_net_1 , \sr_53_[5]_net_1 , \sr_54_[6]_net_1 , 
        \sr_53_[6]_net_1 , \sr_54_[7]_net_1 , \sr_53_[7]_net_1 , 
        \sr_54_[8]_net_1 , \sr_53_[8]_net_1 , \sr_54_[9]_net_1 , 
        \sr_53_[9]_net_1 , \sr_54_[10]_net_1 , \sr_53_[10]_net_1 , 
        \sr_54_[11]_net_1 , \sr_53_[11]_net_1 , \sr_54_[12]_net_1 , 
        \sr_53_[12]_net_1 , \sr_52_[0]_net_1 , \sr_52_[1]_net_1 , 
        \sr_52_[2]_net_1 , \sr_52_[3]_net_1 , \sr_52_[4]_net_1 , 
        \sr_52_[5]_net_1 , \sr_52_[6]_net_1 , \sr_52_[7]_net_1 , 
        \sr_52_[8]_net_1 , \sr_52_[9]_net_1 , \sr_52_[10]_net_1 , 
        \sr_52_[11]_net_1 , \sr_52_[12]_net_1 , \sr_51_[0]_net_1 , 
        \sr_51_[1]_net_1 , \sr_51_[2]_net_1 , \sr_51_[3]_net_1 , 
        \sr_51_[4]_net_1 , \sr_51_[5]_net_1 , \sr_51_[6]_net_1 , 
        \sr_51_[7]_net_1 , \sr_51_[8]_net_1 , \sr_51_[9]_net_1 , 
        \sr_51_[10]_net_1 , \sr_51_[11]_net_1 , \sr_51_[12]_net_1 , 
        \sr_50_[0]_net_1 , \sr_50_[1]_net_1 , \sr_50_[2]_net_1 , 
        \sr_50_[3]_net_1 , \sr_50_[4]_net_1 , \sr_50_[5]_net_1 , 
        \sr_50_[6]_net_1 , \sr_50_[7]_net_1 , \sr_50_[8]_net_1 , 
        \sr_50_[9]_net_1 , \sr_50_[10]_net_1 , \sr_50_[11]_net_1 , 
        \sr_50_[12]_net_1 , \sr_49_[0]_net_1 , \sr_49_[1]_net_1 , 
        \sr_49_[2]_net_1 , \sr_49_[3]_net_1 , \sr_49_[4]_net_1 , 
        \sr_49_[5]_net_1 , \sr_49_[6]_net_1 , \sr_49_[7]_net_1 , 
        \sr_49_[8]_net_1 , \sr_49_[9]_net_1 , \sr_49_[10]_net_1 , 
        \sr_49_[11]_net_1 , \sr_49_[12]_net_1 , \sr_48_[0]_net_1 , 
        \sr_48_[1]_net_1 , \sr_48_[2]_net_1 , \sr_48_[3]_net_1 , 
        \sr_48_[4]_net_1 , \sr_48_[5]_net_1 , \sr_48_[6]_net_1 , 
        \sr_48_[7]_net_1 , \sr_48_[8]_net_1 , \sr_48_[9]_net_1 , 
        \sr_48_[10]_net_1 , \sr_48_[11]_net_1 , \sr_48_[12]_net_1 , 
        \sr_47_[0]_net_1 , \sr_47_[1]_net_1 , \sr_47_[2]_net_1 , 
        \sr_47_[3]_net_1 , \sr_47_[4]_net_1 , \sr_47_[5]_net_1 , 
        \sr_47_[6]_net_1 , \sr_47_[7]_net_1 , \sr_47_[8]_net_1 , 
        \sr_47_[9]_net_1 , \sr_47_[10]_net_1 , \sr_47_[11]_net_1 , 
        \sr_47_[12]_net_1 , \sr_46_[0]_net_1 , \sr_46_[1]_net_1 , 
        \sr_46_[2]_net_1 , \sr_46_[3]_net_1 , \sr_46_[4]_net_1 , 
        \sr_46_[5]_net_1 , \sr_46_[6]_net_1 , \sr_46_[7]_net_1 , 
        \sr_46_[8]_net_1 , \sr_46_[9]_net_1 , \sr_46_[10]_net_1 , 
        \sr_46_[11]_net_1 , \sr_46_[12]_net_1 , \sr_45_[0]_net_1 , 
        \sr_45_[1]_net_1 , \sr_45_[2]_net_1 , \sr_45_[3]_net_1 , 
        \sr_45_[4]_net_1 , \sr_45_[5]_net_1 , \sr_45_[6]_net_1 , 
        \sr_45_[7]_net_1 , \sr_45_[8]_net_1 , \sr_45_[9]_net_1 , 
        \sr_45_[10]_net_1 , \sr_45_[11]_net_1 , \sr_45_[12]_net_1 , 
        \sr_44_[0]_net_1 , \sr_44_[1]_net_1 , \sr_44_[2]_net_1 , 
        \sr_44_[3]_net_1 , \sr_44_[4]_net_1 , \sr_44_[5]_net_1 , 
        \sr_44_[6]_net_1 , \sr_44_[7]_net_1 , \sr_44_[8]_net_1 , 
        \sr_44_[9]_net_1 , \sr_44_[10]_net_1 , \sr_44_[11]_net_1 , 
        \sr_44_[12]_net_1 , \sr_43_[0]_net_1 , \sr_43_[1]_net_1 , 
        \sr_43_[2]_net_1 , \sr_43_[3]_net_1 , \sr_43_[4]_net_1 , 
        \sr_43_[5]_net_1 , \sr_43_[6]_net_1 , \sr_43_[7]_net_1 , 
        \sr_43_[8]_net_1 , \sr_43_[9]_net_1 , \sr_43_[10]_net_1 , 
        \sr_43_[11]_net_1 , \sr_43_[12]_net_1 , \sr_42_[0]_net_1 , 
        \sr_42_[1]_net_1 , \sr_42_[2]_net_1 , \sr_42_[3]_net_1 , 
        \sr_42_[4]_net_1 , \sr_42_[5]_net_1 , \sr_42_[6]_net_1 , 
        \sr_42_[7]_net_1 , \sr_42_[8]_net_1 , \sr_42_[9]_net_1 , 
        \sr_42_[10]_net_1 , \sr_42_[11]_net_1 , \sr_42_[12]_net_1 , 
        \sr_41_[0]_net_1 , \sr_41_[1]_net_1 , \sr_41_[2]_net_1 , 
        \sr_41_[3]_net_1 , \sr_41_[4]_net_1 , \sr_41_[5]_net_1 , 
        \sr_41_[6]_net_1 , \sr_41_[7]_net_1 , \sr_41_[8]_net_1 , 
        \sr_41_[9]_net_1 , \sr_41_[10]_net_1 , \sr_41_[11]_net_1 , 
        \sr_41_[12]_net_1 , \sr_40_[0]_net_1 , \sr_40_[1]_net_1 , 
        \sr_40_[2]_net_1 , \sr_40_[3]_net_1 , \sr_40_[4]_net_1 , 
        \sr_40_[5]_net_1 , \sr_40_[6]_net_1 , \sr_40_[7]_net_1 , 
        \sr_40_[8]_net_1 , \sr_40_[9]_net_1 , \sr_40_[10]_net_1 , 
        \sr_40_[11]_net_1 , \sr_40_[12]_net_1 , \sr_62_[0]_net_1 , 
        \sr_62_[1]_net_1 , \sr_62_[2]_net_1 , \sr_62_[3]_net_1 , 
        \sr_62_[4]_net_1 , \sr_62_[5]_net_1 , \sr_62_[6]_net_1 , 
        \sr_62_[7]_net_1 , \sr_62_[8]_net_1 , \sr_62_[9]_net_1 , 
        \sr_62_[10]_net_1 , \sr_62_[11]_net_1 , \sr_62_[12]_net_1 , 
        \sr_61_[0]_net_1 , \sr_61_[1]_net_1 , \sr_61_[2]_net_1 , 
        \sr_61_[3]_net_1 , \sr_61_[4]_net_1 , \sr_61_[5]_net_1 , 
        \sr_61_[6]_net_1 , \sr_61_[7]_net_1 , \sr_61_[8]_net_1 , 
        \sr_61_[9]_net_1 , \sr_61_[10]_net_1 , \sr_61_[11]_net_1 , 
        \sr_61_[12]_net_1 , \sr_60_[0]_net_1 , \sr_60_[1]_net_1 , 
        \sr_60_[2]_net_1 , \sr_60_[3]_net_1 , \sr_60_[4]_net_1 , 
        \sr_60_[5]_net_1 , \sr_60_[6]_net_1 , \sr_60_[7]_net_1 , 
        \sr_60_[8]_net_1 , \sr_60_[9]_net_1 , \sr_60_[10]_net_1 , 
        \sr_60_[11]_net_1 , \sr_60_[12]_net_1 , \sr_59_[0]_net_1 , 
        \sr_59_[1]_net_1 , \sr_59_[2]_net_1 , \sr_59_[3]_net_1 , 
        \sr_59_[4]_net_1 , \sr_59_[5]_net_1 , \sr_59_[6]_net_1 , 
        \sr_59_[7]_net_1 , \sr_59_[8]_net_1 , \sr_59_[9]_net_1 , 
        \sr_59_[10]_net_1 , \sr_59_[11]_net_1 , \sr_59_[12]_net_1 , 
        \sr_58_[0]_net_1 , \sr_58_[1]_net_1 , \sr_58_[2]_net_1 , 
        \sr_58_[3]_net_1 , \sr_58_[4]_net_1 , \sr_58_[5]_net_1 , 
        \sr_58_[6]_net_1 , \sr_58_[7]_net_1 , \sr_58_[8]_net_1 , 
        \sr_58_[9]_net_1 , \sr_58_[10]_net_1 , \sr_58_[11]_net_1 , 
        \sr_58_[12]_net_1 , \sr_57_[0]_net_1 , \sr_57_[1]_net_1 , 
        \sr_57_[2]_net_1 , \sr_57_[3]_net_1 , \sr_57_[4]_net_1 , 
        \sr_57_[5]_net_1 , \sr_57_[6]_net_1 , \sr_57_[7]_net_1 , 
        \sr_57_[8]_net_1 , \sr_57_[9]_net_1 , \sr_57_[10]_net_1 , 
        \sr_57_[11]_net_1 , \sr_57_[12]_net_1 , \sr_56_[0]_net_1 , 
        \sr_56_[1]_net_1 , \sr_56_[2]_net_1 , \sr_56_[3]_net_1 , 
        \sr_56_[4]_net_1 , \sr_56_[5]_net_1 , \sr_56_[6]_net_1 , 
        \sr_56_[7]_net_1 , \sr_56_[8]_net_1 , \sr_56_[9]_net_1 , 
        \sr_56_[10]_net_1 , \sr_56_[11]_net_1 , \sr_56_[12]_net_1 , 
        \sr_55_[0]_net_1 , \sr_55_[1]_net_1 , \sr_55_[2]_net_1 , 
        \sr_55_[3]_net_1 , \sr_55_[4]_net_1 , \sr_55_[5]_net_1 , 
        \sr_55_[6]_net_1 , \sr_55_[7]_net_1 , \sr_55_[8]_net_1 , 
        \sr_55_[9]_net_1 , \sr_55_[10]_net_1 , \sr_55_[11]_net_1 , 
        \sr_55_[12]_net_1 , GND, VCC;
    
    DFN1E1C0 \sr_41_[5]  (.D(\sr_40_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[5]_net_1 ));
    DFN1E1C0 \sr_15_[3]  (.D(\sr_14_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[3]_net_1 ));
    DFN1E1C0 \sr_36_[5]  (.D(\sr_35_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[5]_net_1 ));
    DFN1E1C0 \sr_57_[5]  (.D(\sr_56_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[5]_net_1 ));
    DFN1E1C0 \sr_45_[11]  (.D(\sr_44_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[11]_net_1 ));
    DFN1E1C0 \sr_39_[6]  (.D(\sr_38_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[6]_net_1 ));
    DFN1E1C0 \sr_36_[4]  (.D(\sr_35_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[4]_net_1 ));
    DFN1E1C0 \sr_42_[4]  (.D(\sr_41_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[4]_net_1 ));
    DFN1E1C0 \sr_9_[3]  (.D(\sr_8_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[3]_net_1 ));
    DFN1E1C0 \sr_6_[4]  (.D(\sr_5_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[4]_net_1 ));
    DFN1E1C0 \sr_32_[3]  (.D(\sr_31_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[3]_net_1 ));
    DFN1E1C0 \sr_52_[6]  (.D(\sr_51_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[6]_net_1 ));
    DFN1E1C0 \sr_21_[9]  (.D(\sr_20_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[9]_net_1 ));
    DFN1E1C0 \sr_47_[12]  (.D(\sr_46_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[12]_net_1 ));
    DFN1E1C0 \sr_22_[4]  (.D(\sr_21_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[4]_net_1 ));
    DFN1E1C0 \sr_10_[1]  (.D(\sr_9_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[1]_net_1 ));
    DFN1E1C0 \sr_5_[4]  (.D(\sr_4_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[4]_net_1 ));
    DFN1E1C0 \sr_62_[6]  (.D(\sr_61_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[6]_net_1 ));
    DFN1E1C0 \sr_58_[2]  (.D(\sr_57_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[2]_net_1 ));
    DFN1E1C0 \sr_55_[0]  (.D(\sr_54_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[0]_net_1 ));
    DFN1E1C0 \sr_27_[3]  (.D(\sr_26_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[3]_net_1 ));
    DFN1E1C0 \sr_21_[1]  (.D(\sr_20_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[1]_net_1 ));
    DFN1E1C0 \sr_37_[9]  (.D(\sr_36_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[9]_net_1 ));
    DFN1E1C0 \sr_48_[10]  (.D(\sr_47_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[10]_net_1 ));
    DFN1E1C0 \sr_60_[5]  (.D(\sr_59_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[5]_net_1 ));
    DFN1E1C0 \sr_30_[5]  (.D(\sr_29_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[5]_net_1 ));
    DFN1E1C0 \sr_14_[4]  (.D(\sr_13_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[4]_net_1 ));
    DFN1E1C0 \sr_24_[8]  (.D(\sr_23_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[8]_net_1 ));
    DFN1E1C0 \sr_30_[4]  (.D(\sr_29_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[4]_net_1 ));
    DFN1E1C0 \sr_37_[6]  (.D(\sr_36_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[6]_net_1 ));
    DFN1E1C0 \sr_42_[6]  (.D(\sr_41_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[6]_net_1 ));
    DFN1E1C0 \sr_58_[4]  (.D(\sr_57_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[4]_net_1 ));
    DFN1E1C0 \sr_57_[10]  (.D(\sr_56_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[10]_net_1 ));
    DFN1E1C0 \sr_43_[7]  (.D(\sr_42_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[7]_net_1 ));
    DFN1E1C0 \sr_44_[2]  (.D(\sr_43_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[2]_net_1 ));
    DFN1E1C0 \sr_53_[7]  (.D(\sr_52_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[7]_net_1 ));
    DFN1E1C0 \sr_59_[1]  (.D(\sr_58_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[1]_net_1 ));
    DFN1E1C0 \sr_27_[10]  (.D(\sr_26_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[10]_net_1 ));
    DFN1E1C0 \sr_53_[8]  (.D(\sr_52_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[8]_net_1 ));
    DFN1E1C0 \sr_16_[4]  (.D(\sr_15_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[4]_net_1 ));
    DFN1E1C0 \sr_10_[11]  (.D(\sr_9_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[11]_net_1 ));
    DFN1E1C0 \sr_26_[8]  (.D(\sr_25_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[8]_net_1 ));
    DFN1E1C0 \sr_63_[7]  (.D(\sr_62_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[7]));
    DFN1E1C0 \sr_28_[7]  (.D(\sr_27_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[7]_net_1 ));
    DFN1E1C0 \sr_63_[8]  (.D(\sr_62_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[8]));
    DFN1E1C0 \sr_24_[0]  (.D(\sr_23_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[0]_net_1 ));
    DFN1E1C0 \sr_46_[2]  (.D(\sr_45_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[2]_net_1 ));
    DFN1E1C0 \sr_13_[5]  (.D(\sr_12_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[5]_net_1 ));
    DFN1E1C0 \sr_0_[2]  (.D(cur_error[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[2]));
    DFN1E1C0 \sr_0_[8]  (.D(cur_error[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[8]));
    DFN1E1C0 \sr_8_[3]  (.D(\sr_7_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[3]_net_1 ));
    DFN1E1C0 \sr_42_[11]  (.D(\sr_41_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[11]_net_1 ));
    DFN1E1C0 \sr_13_[3]  (.D(\sr_12_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[3]_net_1 ));
    DFN1E1C0 \sr_54_[10]  (.D(\sr_53_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[10]_net_1 ));
    DFN1E1C0 \sr_37_[11]  (.D(\sr_36_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[11]_net_1 ));
    DFN1E1C0 \sr_19_[7]  (.D(\sr_18_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[7]_net_1 ));
    DFN1E1C0 \sr_57_[1]  (.D(\sr_56_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[1]_net_1 ));
    DFN1E1C0 \sr_44_[11]  (.D(\sr_43_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[11]_net_1 ));
    DFN1E1C0 \sr_32_[10]  (.D(\sr_31_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[10]_net_1 ));
    DFN1E1C0 \sr_26_[0]  (.D(\sr_25_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[0]_net_1 ));
    DFN1E1C0 \sr_24_[10]  (.D(\sr_23_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[10]_net_1 ));
    DFN1E1C0 \sr_12_[1]  (.D(\sr_11_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[1]_net_1 ));
    DFN1E1C0 \sr_10_[4]  (.D(\sr_9_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[4]_net_1 ));
    DFN1E1C0 \sr_63_[0]  (.D(\sr_62_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[0]));
    DFN1E1C0 \sr_20_[8]  (.D(\sr_19_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[8]_net_1 ));
    DFN1E1C0 \sr_60_[12]  (.D(\sr_59_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[12]_net_1 ));
    DFN1E1C0 \sr_6_[10]  (.D(\sr_5_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[10]_net_1 ));
    DFN1E1C0 \sr_19_[6]  (.D(\sr_18_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[6]_net_1 ));
    DFN1E1C0 \sr_62_[5]  (.D(\sr_61_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[5]_net_1 ));
    DFN1E1C0 \sr_44_[8]  (.D(\sr_43_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[8]_net_1 ));
    DFN1E1C0 \sr_49_[5]  (.D(\sr_48_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[5]_net_1 ));
    DFN1E1C0 \sr_53_[0]  (.D(\sr_52_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[0]_net_1 ));
    DFN1E1C0 \sr_1_[2]  (.D(sr_new[2]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[2]));
    DFN1E1C0 \sr_40_[2]  (.D(\sr_39_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[2]_net_1 ));
    DFN1E1C0 \sr_32_[5]  (.D(\sr_31_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[5]_net_1 ));
    DFN1E1C0 \sr_1_[8]  (.D(sr_new[8]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[8]));
    DFN1E1C0 \sr_18_[12]  (.D(\sr_17_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[12]_net_1 ));
    DFN1E1C0 \sr_60_[10]  (.D(\sr_59_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[10]_net_1 ));
    DFN1E1C0 \sr_32_[4]  (.D(\sr_31_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[4]_net_1 ));
    DFN1E1C0 \sr_54_[3]  (.D(\sr_53_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[3]_net_1 ));
    DFN1E1C0 \sr_29_[9]  (.D(\sr_28_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[9]_net_1 ));
    DFN1E1C0 \sr_24_[2]  (.D(\sr_23_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[2]_net_1 ));
    DFN1E1C0 \sr_18_[9]  (.D(\sr_17_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[9]_net_1 ));
    DFN1E1C0 \sr_7_[9]  (.D(\sr_6_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[9]_net_1 ));
    DFN1E1C0 \sr_63_[10]  (.D(\sr_62_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[10]));
    DFN1E1C0 \sr_24_[5]  (.D(\sr_23_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[5]_net_1 ));
    DFN1E1C0 \sr_46_[8]  (.D(\sr_45_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[8]_net_1 ));
    DFN1E1C0 \sr_59_[11]  (.D(\sr_58_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[11]_net_1 ));
    DFN1E1C0 \sr_17_[7]  (.D(\sr_16_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[7]_net_1 ));
    DFN1E1C0 \sr_14_[8]  (.D(\sr_13_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[8]_net_1 ));
    DFN1E1C0 \sr_41_[3]  (.D(\sr_40_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[3]_net_1 ));
    DFN1E1C0 \sr_20_[0]  (.D(\sr_19_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[0]_net_1 ));
    DFN1E1C0 \sr_48_[0]  (.D(\sr_47_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[0]_net_1 ));
    DFN1E1C0 \sr_29_[1]  (.D(\sr_28_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[1]_net_1 ));
    DFN1E1C0 \sr_3_[10]  (.D(\sr_2_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[10]_net_1 ));
    DFN1E1C0 \sr_29_[11]  (.D(\sr_28_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[11]_net_1 ));
    DFN1E1C0 \sr_35_[1]  (.D(\sr_34_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[1]_net_1 ));
    DFN1E1C0 \sr_17_[6]  (.D(\sr_16_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[6]_net_1 ));
    DFN1E1C0 \sr_2_[3]  (.D(sr_prev[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[3]_net_1 ));
    DFN1E1C0 \sr_56_[3]  (.D(\sr_55_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[3]_net_1 ));
    DFN1E1C0 \sr_47_[5]  (.D(\sr_46_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[5]_net_1 ));
    DFN1E1C0 \sr_35_[2]  (.D(\sr_34_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[2]_net_1 ));
    DFN1E1C0 \sr_35_[12]  (.D(\sr_34_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[12]_net_1 ));
    DFN1E1C0 \sr_26_[2]  (.D(\sr_25_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[2]_net_1 ));
    DFN1E1C0 \sr_6_[2]  (.D(\sr_5_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[2]_net_1 ));
    DFN1E1C0 \sr_6_[8]  (.D(\sr_5_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[8]_net_1 ));
    DFN1E1C0 \sr_35_[7]  (.D(\sr_34_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[7]_net_1 ));
    DFN1E1C0 \sr_26_[5]  (.D(\sr_25_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[5]_net_1 ));
    DFN1E1C0 \sr_16_[8]  (.D(\sr_15_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[8]_net_1 ));
    DFN1E1C0 \sr_52_[12]  (.D(\sr_51_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[12]_net_1 ));
    DFN1E1C0 \sr_5_[2]  (.D(\sr_4_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[2]_net_1 ));
    DFN1E1C0 \sr_5_[8]  (.D(\sr_4_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[8]_net_1 ));
    DFN1E1C0 \sr_27_[9]  (.D(\sr_26_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[9]_net_1 ));
    DFN1E1C0 \sr_18_[11]  (.D(\sr_17_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[11]_net_1 ));
    DFN1E1C0 \sr_3_[9]  (.D(\sr_2_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[9]_net_1 ));
    DFN1E1C0 \sr_2_[11]  (.D(sr_prev[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[11]_net_1 ));
    DFN1E1C0 \sr_40_[8]  (.D(\sr_39_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[8]_net_1 ));
    DFN1E1C0 \sr_22_[12]  (.D(\sr_21_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[12]_net_1 ));
    DFN1E1C0 \sr_45_[9]  (.D(\sr_44_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[9]_net_1 ));
    DFN1E1C0 \sr_2_[12]  (.D(sr_prev[12]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[12]_net_1 ));
    DFN1E1C0 \sr_27_[1]  (.D(\sr_26_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[1]_net_1 ));
    DFN1E1C0 \sr_9_[4]  (.D(\sr_8_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[4]_net_1 ));
    DFN1E1C0 \sr_12_[4]  (.D(\sr_11_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[4]_net_1 ));
    DFN1E1C0 \sr_56_[11]  (.D(\sr_55_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[11]_net_1 ));
    DFN1E1C0 \sr_22_[8]  (.D(\sr_21_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[8]_net_1 ));
    DFN1E1C0 \sr_14_[2]  (.D(\sr_13_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[2]_net_1 ));
    DFN1E1C0 \sr_46_[12]  (.D(\sr_45_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[12]_net_1 ));
    DFN1E1C0 \sr_50_[3]  (.D(\sr_49_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[3]_net_1 ));
    DFN1E1C0 \sr_20_[2]  (.D(\sr_19_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[2]_net_1 ));
    DFN1E1C0 \sr_44_[12]  (.D(\sr_43_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[12]_net_1 ));
    DFN1E1C0 \sr_26_[11]  (.D(\sr_25_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[11]_net_1 ));
    DFN1E1C0 \sr_14_[0]  (.D(\sr_13_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[0]_net_1 ));
    DFN1E1C0 \sr_34_[8]  (.D(\sr_33_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[8]_net_1 ));
    DFN1E1C0 \sr_20_[5]  (.D(\sr_19_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[5]_net_1 ));
    DFN1E1C0 \sr_10_[8]  (.D(\sr_9_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[8]_net_1 ));
    DFN1E1C0 \sr_42_[2]  (.D(\sr_41_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[2]_net_1 ));
    DFN1E1C0 \sr_55_[11]  (.D(\sr_54_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[11]_net_1 ));
    DFN1E1C0 \sr_51_[9]  (.D(\sr_50_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[9]_net_1 ));
    DFN1E1C0 \sr_54_[5]  (.D(\sr_53_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[5]_net_1 ));
    DFN1E1C0 \sr_25_[11]  (.D(\sr_24_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[11]_net_1 ));
    DFN1E1C0 \sr_21_[6]  (.D(\sr_20_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[6]_net_1 ));
    DFN1E1C0 \sr_57_[12]  (.D(\sr_56_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[12]_net_1 ));
    DFN1E1C0 \sr_16_[2]  (.D(\sr_15_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[2]_net_1 ));
    DFN1E1C0 \sr_35_[0]  (.D(\sr_34_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[0]_net_1 ));
    DFN1E1C0 \sr_16_[0]  (.D(\sr_15_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[0]_net_1 ));
    DFN1E1C0 \sr_36_[8]  (.D(\sr_35_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[8]_net_1 ));
    DFN1E1C0 \sr_27_[12]  (.D(\sr_26_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[12]_net_1 ));
    DFN1E1C0 \sr_22_[0]  (.D(\sr_21_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[0]_net_1 ));
    DFN1E1C0 \sr_0__0[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_new_0_0));
    DFN1E1C0 \sr_13_[11]  (.D(\sr_12_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[11]_net_1 ));
    DFN1E1C0 \sr_58_[10]  (.D(\sr_57_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[10]_net_1 ));
    DFN1E1C0 \sr_7_[12]  (.D(\sr_6_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[12]_net_1 ));
    DFN1E1C0 \sr_24_[3]  (.D(\sr_23_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[3]_net_1 ));
    DFN1E1C0 \sr_34_[9]  (.D(\sr_33_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[9]_net_1 ));
    DFN1E1C0 \sr_28_[10]  (.D(\sr_27_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[10]_net_1 ));
    DFN1E1C0 \sr_56_[5]  (.D(\sr_55_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[5]_net_1 ));
    DFN1E1C0 \sr_7_[10]  (.D(\sr_6_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[10]_net_1 ));
    DFN1E1C0 \sr_33_[1]  (.D(\sr_32_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[1]_net_1 ));
    DFN1E1C0 \sr_33_[2]  (.D(\sr_32_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[2]_net_1 ));
    DFN1E1C0 \sr_48_[7]  (.D(\sr_47_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[7]_net_1 ));
    DFN1E1C0 \sr_58_[7]  (.D(\sr_57_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[7]_net_1 ));
    DFN1E1C0 \sr_34_[6]  (.D(\sr_33_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[6]_net_1 ));
    DFN1E1C0 \sr_33_[7]  (.D(\sr_32_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[7]_net_1 ));
    DFN1E1C0 \sr_10_[2]  (.D(\sr_9_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[2]_net_1 ));
    DFN1E1C0 \sr_26_[3]  (.D(\sr_25_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[3]_net_1 ));
    DFN1E1C0 \sr_36_[9]  (.D(\sr_35_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[9]_net_1 ));
    DFN1E1C0 \sr_58_[8]  (.D(\sr_57_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[8]_net_1 ));
    DFN1E1C0 \sr_42_[8]  (.D(\sr_41_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[8]_net_1 ));
    DFN1E1C0 \sr_49_[3]  (.D(\sr_48_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[3]_net_1 ));
    DFN1E1C0 \sr_10_[0]  (.D(\sr_9_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[0]_net_1 ));
    DFN1E1C0 \sr_30_[8]  (.D(\sr_29_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[8]_net_1 ));
    DFN1E1C0 \sr_35_[10]  (.D(\sr_34_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[10]_net_1 ));
    DFN1E1C0 \sr_8_[4]  (.D(\sr_7_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[4]_net_1 ));
    DFN1E1C0 \sr_43_[12]  (.D(\sr_42_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[12]_net_1 ));
    DFN1E1C0 \sr_0_[9]  (.D(cur_error[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[9]));
    DFN1E1C0 \sr_43_[9]  (.D(\sr_42_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[9]_net_1 ));
    DFN1E1C0 \sr_50_[5]  (.D(\sr_49_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[5]_net_1 ));
    DFN1E1C0 \sr_52_[3]  (.D(\sr_51_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[3]_net_1 ));
    DFN1E1C0 \sr_22_[2]  (.D(\sr_21_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[2]_net_1 ));
    DFN1E1C0 \sr_18_[5]  (.D(\sr_17_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[5]_net_1 ));
    DFN1E1C0 \sr_7_[0]  (.D(\sr_6_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[0]_net_1 ));
    DFN1E1C0 \sr_36_[6]  (.D(\sr_35_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[6]_net_1 ));
    DFN1E1C0 \sr_60_[11]  (.D(\sr_59_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[11]_net_1 ));
    DFN1E1C0 \sr_45_[4]  (.D(\sr_44_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[4]_net_1 ));
    DFN1E1C0 \sr_22_[5]  (.D(\sr_21_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[5]_net_1 ));
    DFN1E1C0 \sr_35_[3]  (.D(\sr_34_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[3]_net_1 ));
    DFN1E1C0 \sr_7_[6]  (.D(\sr_6_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[6]_net_1 ));
    DFN1E1C0 \sr_12_[8]  (.D(\sr_11_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[8]_net_1 ));
    DFN1E1C0 \sr_55_[6]  (.D(\sr_54_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[6]_net_1 ));
    DFN1E1C0 \sr_52_[11]  (.D(\sr_51_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[11]_net_1 ));
    DFN1E1C0 \sr_18_[3]  (.D(\sr_17_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[3]_net_1 ));
    DFN1E1C0 \sr_36_[10]  (.D(\sr_35_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[10]_net_1 ));
    DFN1E1C0 \sr_25_[4]  (.D(\sr_24_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[4]_net_1 ));
    DFN1E1C0 \sr_22_[11]  (.D(\sr_21_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[11]_net_1 ));
    DFN1E1C0 \sr_20_[3]  (.D(\sr_19_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[3]_net_1 ));
    DFN1E1C0 \sr_30_[9]  (.D(\sr_29_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[9]_net_1 ));
    DFN1E1C0 \sr_47_[3]  (.D(\sr_46_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[3]_net_1 ));
    DFN1E1C0 \sr_54_[11]  (.D(\sr_53_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[11]_net_1 ));
    DFN1E1C0 \sr_4_[7]  (.D(\sr_3_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[7]_net_1 ));
    DFN1E1C0 \sr_31_[12]  (.D(\sr_30_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[12]_net_1 ));
    DFN1E1C0 \sr_54_[1]  (.D(\sr_53_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[1]_net_1 ));
    DFN1E1C0 \sr_24_[11]  (.D(\sr_23_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[11]_net_1 ));
    DFN1E1C0 \sr_1_[9]  (.D(sr_new[9]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[9]));
    DFN1E1C0 \sr_58_[0]  (.D(\sr_57_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[0]_net_1 ));
    DFN1E1C0 \sr_33_[0]  (.D(\sr_32_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[0]_net_1 ));
    DFN1E1C0 \sr_41_[1]  (.D(\sr_40_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[1]_net_1 ));
    DFN1E1C0 \sr_30_[6]  (.D(\sr_29_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[6]_net_1 ));
    DFN1E1C0 \sr_7_[1]  (.D(\sr_6_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[1]_net_1 ));
    DFN1E1C0 \sr_3_[0]  (.D(\sr_2_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[0]_net_1 ));
    DFN1E1C0 \sr_45_[6]  (.D(\sr_44_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[6]_net_1 ));
    DFN1E1C0 \sr_3_[6]  (.D(\sr_2_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[6]_net_1 ));
    DFN1E1C0 \sr_59_[9]  (.D(\sr_58_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[9]_net_1 ));
    DFN1E1C0 \sr_2_[4]  (.D(sr_prev[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[4]_net_1 ));
    DFN1E1C0 \sr_56_[1]  (.D(\sr_55_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[1]_net_1 ));
    DFN1E1C0 \sr_29_[6]  (.D(\sr_28_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[6]_net_1 ));
    DFN1E1C0 \sr_9_[2]  (.D(\sr_8_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[2]_net_1 ));
    DFN1E1C0 \sr_9_[8]  (.D(\sr_8_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[8]_net_1 ));
    DFN1E1C0 \sr_17_[11]  (.D(\sr_16_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[11]_net_1 ));
    DFN1E1C0 \sr_12_[2]  (.D(\sr_11_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[2]_net_1 ));
    DFN1E1C0 \sr_12_[10]  (.D(\sr_11_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[10]_net_1 ));
    DFN1E1C0 \sr_12_[0]  (.D(\sr_11_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[0]_net_1 ));
    DFN1E1C0 \sr_32_[8]  (.D(\sr_31_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[8]_net_1 ));
    DFN1E1C0 \sr_14_[7]  (.D(\sr_13_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[7]_net_1 ));
    DFN1E1C0 \sr_6_[9]  (.D(\sr_5_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[9]_net_1 ));
    DFN1E1C0 \sr_31_[10]  (.D(\sr_30_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[10]_net_1 ));
    DFN1E1C0 \sr_31_[11]  (.D(\sr_30_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[11]_net_1 ));
    DFN1E1C0 \sr_14_[6]  (.D(\sr_13_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[6]_net_1 ));
    DFN1E1C0 \sr_5_[10]  (.D(\sr_4_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[10]_net_1 ));
    DFN1E1C0 \sr_5_[9]  (.D(\sr_4_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[9]_net_1 ));
    DFN1E1C0 \sr_52_[5]  (.D(\sr_51_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[5]_net_1 ));
    DFN1E1C0 \sr_3_[1]  (.D(\sr_2_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[1]_net_1 ));
    DFN1E1C0 \sr_44_[5]  (.D(\sr_43_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[5]_net_1 ));
    DFN1E1C0 \sr_57_[9]  (.D(\sr_56_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[9]_net_1 ));
    DFN1E1C0 \sr_50_[1]  (.D(\sr_49_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[1]_net_1 ));
    DFN1E1C0 \sr_16_[7]  (.D(\sr_15_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[7]_net_1 ));
    DFN1E1C0 \sr_51_[2]  (.D(\sr_50_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[2]_net_1 ));
    DFN1E1C0 \sr_27_[6]  (.D(\sr_26_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[6]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1C0 \sr_43_[4]  (.D(\sr_42_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[4]_net_1 ));
    DFN1E1C0 \sr_24_[9]  (.D(\sr_23_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[9]_net_1 ));
    DFN1E1C0 \sr_22_[3]  (.D(\sr_21_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[3]_net_1 ));
    DFN1E1C0 \sr_33_[3]  (.D(\sr_32_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[3]_net_1 ));
    DFN1E1C0 \sr_32_[9]  (.D(\sr_31_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[9]_net_1 ));
    DFN1E1C0 \sr_15_[1]  (.D(\sr_14_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[1]_net_1 ));
    DFN1E1C0 \sr_53_[6]  (.D(\sr_52_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[6]_net_1 ));
    DFN1E1C0 \sr_60_[1]  (.D(\sr_59_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[1]_net_1 ));
    DFN1E1C0 \sr_16_[6]  (.D(\sr_15_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[6]_net_1 ));
    DFN1E1C0 \sr_61_[2]  (.D(\sr_60_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[2]_net_1 ));
    DFN1E1C0 \sr_23_[4]  (.D(\sr_22_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[4]_net_1 ));
    DFN1E1C0 \sr_46_[5]  (.D(\sr_45_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[5]_net_1 ));
    DFN1E1C0 \sr_24_[1]  (.D(\sr_23_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[1]_net_1 ));
    DFN1E1C0 \sr_63_[6]  (.D(\sr_62_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[6]));
    DFN1E1C0 \sr_49_[12]  (.D(\sr_48_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[12]_net_1 ));
    DFN1E1C0 \sr_56_[12]  (.D(\sr_55_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[12]_net_1 ));
    DFN1E1C0 \sr_54_[12]  (.D(\sr_53_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[12]_net_1 ));
    DFN1E1C0 \sr_35_[5]  (.D(\sr_34_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[5]_net_1 ));
    DFN1E1C0 \sr_15_[12]  (.D(\sr_14_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[12]_net_1 ));
    DFN1E1C0 \sr_32_[6]  (.D(\sr_31_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[6]_net_1 ));
    DFN1E1C0 \sr_26_[12]  (.D(\sr_25_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[12]_net_1 ));
    DFN1E1C0 \sr_35_[4]  (.D(\sr_34_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[4]_net_1 ));
    DFN1E1C0 \sr_26_[9]  (.D(\sr_25_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[9]_net_1 ));
    DFN1E1C0 \sr_24_[12]  (.D(\sr_23_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[12]_net_1 ));
    DFN1E1C0 \sr_51_[4]  (.D(\sr_50_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[4]_net_1 ));
    DFN1E1C0 \sr_10_[7]  (.D(\sr_9_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[7]_net_1 ));
    DFN1E1C0 \sr_8_[2]  (.D(\sr_7_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[2]_net_1 ));
    DFN1E1C0 \sr_40_[12]  (.D(\sr_39_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[12]_net_1 ));
    DFN1E1C0 \sr_8_[8]  (.D(\sr_7_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[8]_net_1 ));
    DFN1E1C0 \sr_26_[1]  (.D(\sr_25_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[1]_net_1 ));
    DFN1E1C0 \sr_61_[4]  (.D(\sr_60_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[4]_net_1 ));
    DFN1E1C0 \sr_0_[0]  (.D(cur_error[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[0]));
    DFN1E1C0 \sr_43_[6]  (.D(\sr_42_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[6]_net_1 ));
    DFN1E1C0 \sr_10_[6]  (.D(\sr_9_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[6]_net_1 ));
    DFN1E1C0 \sr_21_[7]  (.D(\sr_20_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[7]_net_1 ));
    DFN1E1C0 \sr_0_[6]  (.D(cur_error[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[6]));
    DFN1E1C0 \sr_40_[5]  (.D(\sr_39_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[5]_net_1 ));
    DFN1E1C0 \sr_40_[10]  (.D(\sr_39_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[10]_net_1 ));
    DFN1E1C0 \sr_43_[10]  (.D(\sr_42_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[10]_net_1 ));
    DFN1E1C0 \sr_38_[1]  (.D(\sr_37_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[1]_net_1 ));
    DFN1E1C0 \sr_49_[1]  (.D(\sr_48_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[1]_net_1 ));
    DFN1E1C0 \sr_63_[11]  (.D(\sr_62_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[11]));
    DFN1E1C0 \sr_20_[9]  (.D(\sr_19_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[9]_net_1 ));
    DFN1E1C0 \sr_38_[2]  (.D(\sr_37_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[2]_net_1 ));
    DFN1E1C0 \sr_38_[7]  (.D(\sr_37_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[7]_net_1 ));
    DFN1E1C0 \sr_52_[1]  (.D(\sr_51_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[1]_net_1 ));
    DFN1E1C0 \sr_20_[1]  (.D(\sr_19_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[1]_net_1 ));
    DFN1E1C0 \sr_1_[0]  (.D(sr_new[0]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[0]));
    DFN1E1C0 \sr_61_[9]  (.D(\sr_60_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[9]_net_1 ));
    DFN1E1C0 \sr_0_[1]  (.D(cur_error[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[1]));
    DFN1E1C0 \sr_15_[4]  (.D(\sr_14_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[4]_net_1 ));
    DFN1E1C0 \sr_1_[6]  (.D(sr_new[6]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[6]));
    DFN1E1C0 \sr_62_[1]  (.D(\sr_61_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[1]_net_1 ));
    DFN1E1C0 \sr_25_[8]  (.D(\sr_24_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[8]_net_1 ));
    DFN1E1C0 \sr_48_[9]  (.D(\sr_47_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[9]_net_1 ));
    DFN1E1C0 \sr_1_[11]  (.D(sr_new[11]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_prev[11]));
    DFN1E1C0 \sr_49_[10]  (.D(\sr_48_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[10]_net_1 ));
    DFN1E1C0 \sr_53_[12]  (.D(\sr_52_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[12]_net_1 ));
    DFN1E1C0 \sr_13_[1]  (.D(\sr_12_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[1]_net_1 ));
    DFN1E1C0 \sr_7_[5]  (.D(\sr_6_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[5]_net_1 ));
    DFN1E1C0 \sr_5_[12]  (.D(\sr_4_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[12]_net_1 ));
    DFN1E1C0 \sr_47_[1]  (.D(\sr_46_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[1]_net_1 ));
    DFN1E1C0 \sr_23_[12]  (.D(\sr_22_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[12]_net_1 ));
    DFN1E1C0 \sr_63_[5]  (.D(\sr_62_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[5]));
    DFN1E1C0 \sr_45_[2]  (.D(\sr_44_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[2]_net_1 ));
    DFN1E1C0 \sr_2_[2]  (.D(sr_prev[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[2]_net_1 ));
    DFN1E1C0 \sr_2_[8]  (.D(sr_prev[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[8]_net_1 ));
    DFN1E1C0 \sr_11_[9]  (.D(\sr_10_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[9]_net_1 ));
    DFN1E1C0 \sr_33_[5]  (.D(\sr_32_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[5]_net_1 ));
    DFN1E1C0 \sr_59_[2]  (.D(\sr_58_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[2]_net_1 ));
    DFN1E1C0 \sr_12_[7]  (.D(\sr_11_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[7]_net_1 ));
    DFN1E1C0 \sr_6_[0]  (.D(\sr_5_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[0]_net_1 ));
    DFN1E1C0 \sr_41_[0]  (.D(\sr_40_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[0]_net_1 ));
    DFN1E1C0 \sr_1_[1]  (.D(sr_new[1]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[1]));
    DFN1E1C0 \sr_33_[4]  (.D(\sr_32_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[4]_net_1 ));
    DFN1E1C0 \sr_9_[12]  (.D(\sr_8_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[12]_net_1 ));
    DFN1E1C0 \sr_25_[0]  (.D(\sr_24_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[0]_net_1 ));
    DFN1E1C0 \sr_6_[6]  (.D(\sr_5_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[6]_net_1 ));
    DFN1E1C0 \sr_15_[10]  (.D(\sr_14_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[10]_net_1 ));
    DFN1E1C0 \sr_12_[6]  (.D(\sr_11_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[6]_net_1 ));
    DFN1E1C0 \sr_61_[3]  (.D(\sr_60_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[3]_net_1 ));
    DFN1E1C0 \sr_5_[0]  (.D(\sr_4_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[0]_net_1 ));
    DFN1E1C0 \sr_44_[3]  (.D(\sr_43_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[3]_net_1 ));
    DFN1E1C0 \sr_38_[0]  (.D(\sr_37_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[0]_net_1 ));
    DFN1E1C0 \sr_42_[5]  (.D(\sr_41_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[5]_net_1 ));
    DFN1E1C0 \sr_5_[6]  (.D(\sr_4_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[6]_net_1 ));
    DFN1E1C0 \sr_3_[5]  (.D(\sr_2_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[5]_net_1 ));
    DFN1E1C0 \sr_4_[3]  (.D(\sr_3_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[3]_net_1 ));
    DFN1E1C0 \sr_9_[9]  (.D(\sr_8_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[9]_net_1 ));
    DFN1E1C0 \sr_37_[10]  (.D(\sr_36_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[10]_net_1 ));
    DFN1E1C0 \sr_22_[9]  (.D(\sr_21_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[9]_net_1 ));
    DFN1E1C0 \sr_59_[4]  (.D(\sr_58_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[4]_net_1 ));
    DFN1E1C0 \sr_16_[10]  (.D(\sr_15_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[10]_net_1 ));
    DFN1E1C0 \sr_57_[2]  (.D(\sr_56_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[2]_net_1 ));
    DFN1E1C0 \sr_46_[3]  (.D(\sr_45_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[3]_net_1 ));
    DFN1E1C0 \sr_6_[1]  (.D(\sr_5_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[1]_net_1 ));
    DFN1E1C0 \sr_45_[8]  (.D(\sr_44_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[8]_net_1 ));
    DFN1E1C0 \sr_22_[1]  (.D(\sr_21_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[1]_net_1 ));
    DFN1E1C0 \sr_29_[7]  (.D(\sr_28_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[7]_net_1 ));
    DFN1E1C0 \sr_11_[12]  (.D(\sr_10_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[12]_net_1 ));
    DFN1E1C0 \sr_5_[1]  (.D(\sr_4_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[1]_net_1 ));
    DFN1E1C0 \sr_4_[10]  (.D(\sr_3_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[10]_net_1 ));
    DFN1E1C0 \sr_55_[3]  (.D(\sr_54_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[3]_net_1 ));
    DFN1E1C0 \sr_25_[2]  (.D(\sr_24_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[2]_net_1 ));
    DFN1E1C0 \sr_13_[4]  (.D(\sr_12_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[4]_net_1 ));
    DFN1E1C0 \sr_62_[10]  (.D(\sr_61_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[10]_net_1 ));
    DFN1E1C0 \sr_23_[8]  (.D(\sr_22_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[8]_net_1 ));
    DFN1E1C0 \sr_25_[5]  (.D(\sr_24_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[5]_net_1 ));
    DFN1E1C0 \sr_15_[8]  (.D(\sr_14_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[8]_net_1 ));
    DFN1E1C0 \sr_34_[10]  (.D(\sr_33_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[10]_net_1 ));
    DFN1E1C0 \sr_57_[4]  (.D(\sr_56_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[4]_net_1 ));
    DFN1E1C0 \sr_40_[3]  (.D(\sr_39_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[3]_net_1 ));
    DFN1E1C0 \sr_48_[4]  (.D(\sr_47_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[4]_net_1 ));
    DFN1E1C0 \sr_38_[3]  (.D(\sr_37_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[3]_net_1 ));
    DFN1E1C0 \sr_43_[2]  (.D(\sr_42_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[2]_net_1 ));
    DFN1E1C0 \sr_58_[6]  (.D(\sr_57_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[6]_net_1 ));
    DFN1E1C0 \sr_54_[9]  (.D(\sr_53_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[9]_net_1 ));
    DFN1E1C0 \sr_28_[4]  (.D(\sr_27_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[4]_net_1 ));
    DFN1E1C0 \sr_27_[7]  (.D(\sr_26_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[7]_net_1 ));
    DFN1E1C0 \sr_24_[6]  (.D(\sr_23_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[6]_net_1 ));
    DFN1E1C0 \sr_40_[11]  (.D(\sr_39_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[11]_net_1 ));
    DFN1E1C0 \sr_11_[10]  (.D(\sr_10_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[10]_net_1 ));
    DFN1E1C0 \sr_23_[0]  (.D(\sr_22_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[0]_net_1 ));
    DFN1E1C0 \sr_11_[11]  (.D(\sr_10_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[11]_net_1 ));
    DFN1E1C0 \sr_59_[12]  (.D(\sr_58_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[12]_net_1 ));
    DFN1E1C0 \sr_8_[9]  (.D(\sr_7_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[9]_net_1 ));
    DFN1E1C0 \sr_1_[10]  (.D(sr_new[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_prev[10]));
    DFN1E1C0 \sr_41_[7]  (.D(\sr_40_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[7]_net_1 ));
    DFN1E1C0 \sr_29_[12]  (.D(\sr_28_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[12]_net_1 ));
    DFN1E1C0 \sr_19_[9]  (.D(\sr_18_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[9]_net_1 ));
    DFN1E1C0 \sr_56_[9]  (.D(\sr_55_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[9]_net_1 ));
    DFN1E1C0 \sr_51_[7]  (.D(\sr_50_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[7]_net_1 ));
    DFN1E1C0 \sr_39_[11]  (.D(\sr_38_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[11]_net_1 ));
    DFN1E1C0 \sr_26_[6]  (.D(\sr_25_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[6]_net_1 ));
    DFN1E1C0 \sr_51_[8]  (.D(\sr_50_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[8]_net_1 ));
    DFN1E1C0 \sr_50_[12]  (.D(\sr_49_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[12]_net_1 ));
    DFN1E1C0 \sr_49_[0]  (.D(\sr_48_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[0]_net_1 ));
    DFN1E1C0 \sr_0_[5]  (.D(cur_error[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[5]));
    DFN1E1C0 \sr_15_[2]  (.D(\sr_14_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[2]_net_1 ));
    DFN1E1C0 \sr_61_[7]  (.D(\sr_60_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[7]_net_1 ));
    DFN1E1C0 \sr_48_[6]  (.D(\sr_47_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[6]_net_1 ));
    DFN1E1C0 \sr_15_[0]  (.D(\sr_14_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[0]_net_1 ));
    DFN1E1C0 \sr_35_[8]  (.D(\sr_34_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[8]_net_1 ));
    DFN1E1C0 \sr_61_[8]  (.D(\sr_60_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[8]_net_1 ));
    DFN1E1C0 \sr_20_[12]  (.D(\sr_19_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[12]_net_1 ));
    DFN1E1C0 \sr_43_[8]  (.D(\sr_42_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[8]_net_1 ));
    DFN1E1C0 \sr_11_[5]  (.D(\sr_10_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[5]_net_1 ));
    DFN1E1C0 \sr_50_[10]  (.D(\sr_49_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[10]_net_1 ));
    DFN1E1C0 \sr_55_[5]  (.D(\sr_54_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[5]_net_1 ));
    DFN1E1C0 \sr_53_[10]  (.D(\sr_52_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[10]_net_1 ));
    DFN1E1C0 \sr_48_[12]  (.D(\sr_47_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[12]_net_1 ));
    DFN1E1C0 \sr_32_[12]  (.D(\sr_31_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[12]_net_1 ));
    DFN1E1C0 \sr_11_[3]  (.D(\sr_10_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[3]_net_1 ));
    DFN1E1C0 \sr_0_[11]  (.D(cur_error[11]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable), .Q(sr_new[11]));
    DFN1E1C0 \sr_20_[10]  (.D(\sr_19_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[10]_net_1 ));
    DFN1E1C0 \sr_50_[9]  (.D(\sr_49_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[9]_net_1 ));
    DFN1E1C0 \sr_17_[9]  (.D(\sr_16_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[9]_net_1 ));
    DFN1E1C0 \sr_23_[10]  (.D(\sr_22_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[10]_net_1 ));
    DFN1E1C0 \sr_20_[6]  (.D(\sr_19_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[6]_net_1 ));
    DFN1E1C0 \sr_53_[3]  (.D(\sr_52_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[3]_net_1 ));
    DFN1E1C0 \sr_23_[2]  (.D(\sr_22_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[2]_net_1 ));
    DFN1E1C0 \sr_1_[5]  (.D(sr_new[5]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[5]));
    DFN1E1C0 \sr_61_[0]  (.D(\sr_60_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[0]_net_1 ));
    DFN1E1C0 \sr_47_[0]  (.D(\sr_46_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[0]_net_1 ));
    DFN1E1C0 \sr_23_[5]  (.D(\sr_22_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[5]_net_1 ));
    DFN1E1C0 \sr_42_[3]  (.D(\sr_41_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[3]_net_1 ));
    DFN1E1C0 \sr_25_[3]  (.D(\sr_24_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[3]_net_1 ));
    DFN1E1C0 \sr_35_[9]  (.D(\sr_34_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[9]_net_1 ));
    DFN1E1C0 \sr_13_[8]  (.D(\sr_12_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[8]_net_1 ));
    DFN1E1C0 \sr_36_[11]  (.D(\sr_35_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[11]_net_1 ));
    DFN1E1C0 \sr_51_[0]  (.D(\sr_50_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[0]_net_1 ));
    DFN1E1C0 \sr_18_[1]  (.D(\sr_17_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[1]_net_1 ));
    DFN1E1C0 \sr_2_[9]  (.D(sr_prev[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[9]_net_1 ));
    DFN1E1C0 \sr_9_[0]  (.D(\sr_8_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[0]_net_1 ));
    DFN1E1C0 \sr_59_[10]  (.D(\sr_58_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[10]_net_1 ));
    DFN1E1C0 \sr_35_[11]  (.D(\sr_34_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[11]_net_1 ));
    DFN1E1C0 \sr_35_[6]  (.D(\sr_34_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_35_[6]_net_1 ));
    DFN1E1C0 \sr_9_[6]  (.D(\sr_8_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[6]_net_1 ));
    DFN1E1C0 \sr_29_[10]  (.D(\sr_28_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[10]_net_1 ));
    DFN1E1C0 \sr_44_[1]  (.D(\sr_43_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[1]_net_1 ));
    DFN1E1C0 \sr_38_[5]  (.D(\sr_37_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[5]_net_1 ));
    DFN1E1C0 \sr_37_[12]  (.D(\sr_36_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[12]_net_1 ));
    DFN1E1C0 \sr_6_[5]  (.D(\sr_5_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[5]_net_1 ));
    DFN1E1C0 \sr_48_[11]  (.D(\sr_47_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[11]_net_1 ));
    DFN1E1C0 \sr_38_[4]  (.D(\sr_37_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[4]_net_1 ));
    DFN1E1C0 \sr_4_[4]  (.D(\sr_3_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[4]_net_1 ));
    DFN1E1C0 \sr_38_[10]  (.D(\sr_37_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[10]_net_1 ));
    DFN1E1C0 \sr_5_[5]  (.D(\sr_4_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[5]_net_1 ));
    DFN1E1C0 \sr_13_[2]  (.D(\sr_12_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[2]_net_1 ));
    DFN1E1C0 \sr_46_[1]  (.D(\sr_45_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[1]_net_1 ));
    DFN1E1C0 \sr_9_[1]  (.D(\sr_8_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[1]_net_1 ));
    DFN1E1C0 \sr_13_[0]  (.D(\sr_12_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[0]_net_1 ));
    DFN1E1C0 \sr_33_[8]  (.D(\sr_32_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[8]_net_1 ));
    DFN1E1C0 \sr_49_[7]  (.D(\sr_48_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[7]_net_1 ));
    DFN1E1C0 \sr_59_[7]  (.D(\sr_58_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[7]_net_1 ));
    DFN1E1C0 \sr_52_[9]  (.D(\sr_51_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[9]_net_1 ));
    DFN1E1C0 \sr_59_[8]  (.D(\sr_58_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[8]_net_1 ));
    DFN1E1C0 \sr_53_[5]  (.D(\sr_52_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[5]_net_1 ));
    DFN1E1C0 \sr_22_[6]  (.D(\sr_21_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[6]_net_1 ));
    DFN1E1C0 \sr_55_[1]  (.D(\sr_54_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[1]_net_1 ));
    DFN1E1C0 \sr_54_[2]  (.D(\sr_53_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[2]_net_1 ));
    DFN1E1C0 \sr_43_[11]  (.D(\sr_42_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[11]_net_1 ));
    DFN1E1C0 \sr_8_[0]  (.D(\sr_7_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[0]_net_1 ));
    DFN1E1C0 \sr_23_[3]  (.D(\sr_22_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[3]_net_1 ));
    DFN1E1C0 \sr_40_[1]  (.D(\sr_39_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[1]_net_1 ));
    DFN1E1C0 \sr_33_[9]  (.D(\sr_32_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[9]_net_1 ));
    DFN1E1C0 \sr_19_[5]  (.D(\sr_18_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[5]_net_1 ));
    DFN1E1C0 \sr_18_[4]  (.D(\sr_17_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[4]_net_1 ));
    DFN1E1C0 \sr_28_[8]  (.D(\sr_27_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[8]_net_1 ));
    DFN1E1C0 \sr_8_[6]  (.D(\sr_7_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[6]_net_1 ));
    DFN1E1C0 \sr_32_[11]  (.D(\sr_31_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[11]_net_1 ));
    DFN1E1C0 \sr_61_[12]  (.D(\sr_60_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[12]_net_1 ));
    DFN1E1C0 \sr_19_[3]  (.D(\sr_18_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[3]_net_1 ));
    DFN1E1C0 \sr_8_[11]  (.D(\sr_7_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[11]_net_1 ));
    DFN1E1C0 \sr_47_[7]  (.D(\sr_46_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[7]_net_1 ));
    DFN1E1C0 \sr_57_[7]  (.D(\sr_56_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[7]_net_1 ));
    DFN1E1C0 \sr_56_[2]  (.D(\sr_55_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[2]_net_1 ));
    DFN1E1C0 \sr_17_[10]  (.D(\sr_16_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[10]_net_1 ));
    DFN1E1C0 \sr_57_[8]  (.D(\sr_56_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[8]_net_1 ));
    DFN1E1C0 \sr_48_[2]  (.D(\sr_47_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[2]_net_1 ));
    DFN1E1C0 \sr_15_[7]  (.D(\sr_14_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[7]_net_1 ));
    DFN1E1C0 \sr_34_[11]  (.D(\sr_33_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[11]_net_1 ));
    DFN1E1C0 \sr_33_[6]  (.D(\sr_32_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[6]_net_1 ));
    DFN1E1C0 \sr_54_[4]  (.D(\sr_53_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[4]_net_1 ));
    DFN1E1C0 \sr_15_[6]  (.D(\sr_14_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[6]_net_1 ));
    DFN1E1C0 \sr_59_[0]  (.D(\sr_58_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[0]_net_1 ));
    DFN1E1C0 \sr_50_[11]  (.D(\sr_49_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[11]_net_1 ));
    DFN1E1C0 \sr_45_[5]  (.D(\sr_44_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[5]_net_1 ));
    DFN1E1C0 \sr_8_[1]  (.D(\sr_7_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[1]_net_1 ));
    DFN1E1C0 \sr_31_[1]  (.D(\sr_30_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[1]_net_1 ));
    DFN1E1C0 \sr_28_[0]  (.D(\sr_27_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[0]_net_1 ));
    DFN1E1C0 \sr_17_[5]  (.D(\sr_16_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[5]_net_1 ));
    DFN1E1C0 \sr_24_[7]  (.D(\sr_23_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[7]_net_1 ));
    DFN1E1C0 \sr_20_[11]  (.D(\sr_19_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[11]_net_1 ));
    DFN1E1C0 \sr_31_[2]  (.D(\sr_30_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[2]_net_1 ));
    DFN1E1C0 \sr_17_[3]  (.D(\sr_16_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[3]_net_1 ));
    DFN1E1C0 \sr_56_[4]  (.D(\sr_55_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[4]_net_1 ));
    DFN1E1C0 \sr_31_[7]  (.D(\sr_30_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[7]_net_1 ));
    DFN1E1C0 \sr_25_[9]  (.D(\sr_24_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[9]_net_1 ));
    DFN1E1C0 \sr_61_[10]  (.D(\sr_60_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[10]_net_1 ));
    DFN1E1C0 \sr_50_[2]  (.D(\sr_49_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[2]_net_1 ));
    DFN1E1C0 \sr_14_[10]  (.D(\sr_13_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[10]_net_1 ));
    DFN1E1C0 \sr_61_[11]  (.D(\sr_60_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[11]_net_1 ));
    DFN1E1C0 \sr_25_[1]  (.D(\sr_24_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[1]_net_1 ));
    DFN1E1C0 \sr_60_[2]  (.D(\sr_59_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[2]_net_1 ));
    DFN1E1C0 \sr_26_[7]  (.D(\sr_25_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[7]_net_1 ));
    DFN1E1C0 \sr_2_[0]  (.D(sr_prev[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[0]_net_1 ));
    DFN1E1C0 \sr_41_[9]  (.D(\sr_40_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[9]_net_1 ));
    DFN1E1C0 \sr_57_[0]  (.D(\sr_56_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[0]_net_1 ));
    DFN1E1C0 \sr_48_[8]  (.D(\sr_47_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[8]_net_1 ));
    DFN1E1C0 \sr_53_[1]  (.D(\sr_52_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[1]_net_1 ));
    DFN1E1C0 \sr_2_[6]  (.D(sr_prev[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[6]_net_1 ));
    DFN1E1C0 \sr_7_[7]  (.D(\sr_6_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[7]_net_1 ));
    DFN1E1C0 \sr_42_[1]  (.D(\sr_41_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[1]_net_1 ));
    DFN1E1C0 \sr_63_[1]  (.D(\sr_62_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[1]));
    DFN1E1C0 \sr_50_[4]  (.D(\sr_49_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[4]_net_1 ));
    DFN1E1C0 \sr_58_[12]  (.D(\sr_57_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[12]_net_1 ));
    DFN1E1C0 \sr_58_[3]  (.D(\sr_57_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[3]_net_1 ));
    DFN1E1C0 \sr_28_[2]  (.D(\sr_27_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[2]_net_1 ));
    DFN1E1C0 \sr_4_[2]  (.D(\sr_3_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[2]_net_1 ));
    DFN1E1C0 \sr_4_[8]  (.D(\sr_3_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[8]_net_1 ));
    DFN1E1C0 \sr_28_[5]  (.D(\sr_27_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[5]_net_1 ));
    DFN1E1C0 \sr_28_[12]  (.D(\sr_27_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[12]_net_1 ));
    DFN1E1C0 \sr_60_[4]  (.D(\sr_59_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[4]_net_1 ));
    DFN1E1C0 \sr_19_[11]  (.D(\sr_18_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[11]_net_1 ));
    DFN1E1C0 \sr_14_[9]  (.D(\sr_13_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[9]_net_1 ));
    DFN1E1C0 \sr_18_[8]  (.D(\sr_17_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[8]_net_1 ));
    DFN1E1C0 \sr_47_[11]  (.D(\sr_46_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[11]_net_1 ));
    DFN1E1C0 \sr_20_[7]  (.D(\sr_19_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[7]_net_1 ));
    DFN1E1C0 \sr_2_[1]  (.D(sr_prev[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[1]_net_1 ));
    DFN1E1C0 \sr_31_[0]  (.D(\sr_30_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[0]_net_1 ));
    DFN1E1C0 \sr_42_[10]  (.D(\sr_41_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[10]_net_1 ));
    DFN1E1C0 \sr_44_[0]  (.D(\sr_43_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[0]_net_1 ));
    DFN1E1C0 \sr_13_[7]  (.D(\sr_12_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[7]_net_1 ));
    DFN1E1C0 \sr_36_[12]  (.D(\sr_35_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[12]_net_1 ));
    DFN1E1C0 \sr_9_[5]  (.D(\sr_8_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[5]_net_1 ));
    DFN1E1C0 \sr_34_[12]  (.D(\sr_33_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[12]_net_1 ));
    DFN1E1C0 \sr_3_[7]  (.D(\sr_2_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[7]_net_1 ));
    DFN1E1C0 \sr_13_[6]  (.D(\sr_12_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[6]_net_1 ));
    DFN1E1C0 \sr_16_[9]  (.D(\sr_15_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[9]_net_1 ));
    DFN1E1C0 \sr_12_[12]  (.D(\sr_11_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[12]_net_1 ));
    DFN1E1C0 \sr_43_[5]  (.D(\sr_42_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[5]_net_1 ));
    DFN1E1C0 \sr_46_[0]  (.D(\sr_45_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[0]_net_1 ));
    DFN1E1C0 \sr_52_[2]  (.D(\sr_51_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[2]_net_1 ));
    DFN1E1C0 \sr_60_[9]  (.D(\sr_59_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[9]_net_1 ));
    DFN1E1C0 \sr_4_[12]  (.D(\sr_3_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[12]_net_1 ));
    DFN1E1C0 \sr_58_[11]  (.D(\sr_57_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[11]_net_1 ));
    DFN1E1C0 \sr_3_[12]  (.D(\sr_2_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[12]_net_1 ));
    DFN1E1C0 \sr_23_[9]  (.D(\sr_22_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[9]_net_1 ));
    DFN1E1C0 \sr_28_[11]  (.D(\sr_27_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[11]_net_1 ));
    DFN1E1C0 \sr_62_[2]  (.D(\sr_61_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[2]_net_1 ));
    DFN1E1C0 \sr_16_[11]  (.D(\sr_15_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[11]_net_1 ));
    DFN1E1C0 \sr_1_[12]  (.D(sr_new_0_0), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_prev[12]));
    DFN1E1C0 \sr_18_[2]  (.D(\sr_17_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[2]_net_1 ));
    DFN1E1C0 \sr_39_[1]  (.D(\sr_38_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[1]_net_1 ));
    DFN1E1C0 \sr_23_[1]  (.D(\sr_22_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[1]_net_1 ));
    DFN1E1C0 \sr_18_[0]  (.D(\sr_17_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[0]_net_1 ));
    DFN1E1C0 \sr_38_[8]  (.D(\sr_37_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[8]_net_1 ));
    DFN1E1C0 \sr_8_[10]  (.D(\sr_7_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[10]_net_1 ));
    DFN1E1C0 \sr_10_[9]  (.D(\sr_9_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[9]_net_1 ));
    DFN1E1C0 \sr_45_[12]  (.D(\sr_44_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[12]_net_1 ));
    DFN1E1C0 \sr_39_[2]  (.D(\sr_38_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[2]_net_1 ));
    DFN1E1C0 \sr_8_[12]  (.D(\sr_7_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[12]_net_1 ));
    DFN1E1C0 \sr_15_[11]  (.D(\sr_14_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[11]_net_1 ));
    DFN1E1C0 \sr_39_[7]  (.D(\sr_38_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[7]_net_1 ));
    DFN1E1C0 \sr_52_[4]  (.D(\sr_51_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[4]_net_1 ));
    DFN1E1C0 \sr_41_[4]  (.D(\sr_40_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[4]_net_1 ));
    DFN1E1C0 \sr_58_[5]  (.D(\sr_57_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[5]_net_1 ));
    DFN1E1C0 \sr_40_[0]  (.D(\sr_39_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[0]_net_1 ));
    DFN1E1C0 \sr_31_[3]  (.D(\sr_30_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[3]_net_1 ));
    DFN1E1C0 \sr_51_[6]  (.D(\sr_50_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[6]_net_1 ));
    DFN1E1C0 \sr_17_[12]  (.D(\sr_16_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[12]_net_1 ));
    DFN1E1C0 \sr_45_[3]  (.D(\sr_44_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[3]_net_1 ));
    DFN1E1C0 \sr_62_[4]  (.D(\sr_61_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[4]_net_1 ));
    DFN1E1C0 \sr_21_[4]  (.D(\sr_20_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[4]_net_1 ));
    DFN1E1C0 \sr_60_[3]  (.D(\sr_59_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[3]_net_1 ));
    DFN1E1C0 \sr_22_[7]  (.D(\sr_21_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[7]_net_1 ));
    DFN1E1C0 \sr_61_[6]  (.D(\sr_60_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[6]_net_1 ));
    DFN1E1C0 \sr_49_[9]  (.D(\sr_48_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[9]_net_1 ));
    DFN1E1C0 \sr_18_[10]  (.D(\sr_17_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[10]_net_1 ));
    DFN1E1C0 \sr_8_[5]  (.D(\sr_7_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[5]_net_1 ));
    DFN1E1C0 \sr_33_[12]  (.D(\sr_32_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[12]_net_1 ));
    DFN1E1C0 \sr_28_[3]  (.D(\sr_27_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[3]_net_1 ));
    DFN1E1C0 \sr_38_[9]  (.D(\sr_37_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[9]_net_1 ));
    DFN1E1C0 \sr_53_[11]  (.D(\sr_52_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[11]_net_1 ));
    DFN1E1C0 \sr_37_[1]  (.D(\sr_36_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[1]_net_1 ));
    DFN1E1C0 \sr_37_[2]  (.D(\sr_36_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[2]_net_1 ));
    DFN1E1C0 \sr_23_[11]  (.D(\sr_22_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[11]_net_1 ));
    DFN1E1C0 \sr_3_[11]  (.D(\sr_2_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[11]_net_1 ));
    DFN1E1C0 \sr_37_[7]  (.D(\sr_36_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[7]_net_1 ));
    DFN1E1C0 \sr_38_[6]  (.D(\sr_37_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[6]_net_1 ));
    DFN1E1C0 \sr_41_[6]  (.D(\sr_40_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[6]_net_1 ));
    DFN1E1C0 \sr_44_[7]  (.D(\sr_43_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[7]_net_1 ));
    DFN1E1C0 \sr_54_[7]  (.D(\sr_53_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[7]_net_1 ));
    DFN1E1C0 \sr_0_[7]  (.D(cur_error[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[7]));
    DFN1E1C0 \sr_9_[11]  (.D(\sr_8_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[11]_net_1 ));
    DFN1E1C0 \sr_62_[9]  (.D(\sr_61_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[9]_net_1 ));
    DFN1E1C0 \sr_54_[8]  (.D(\sr_53_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[8]_net_1 ));
    DFN1E1C0 \sr_39_[0]  (.D(\sr_38_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[0]_net_1 ));
    DFN1E1C0 \sr_47_[9]  (.D(\sr_46_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[9]_net_1 ));
    DFN1E1C0 \sr_6_[12]  (.D(\sr_5_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[12]_net_1 ));
    DFN1E1C0 \sr_7_[11]  (.D(\sr_6_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[11]_net_1 ));
    DFN1E1C0 \sr_46_[7]  (.D(\sr_45_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[7]_net_1 ));
    DFN1E1C0 \sr_14_[5]  (.D(\sr_13_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[5]_net_1 ));
    DFN1E1C0 \sr_56_[7]  (.D(\sr_55_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[7]_net_1 ));
    DFN1E1C0 \sr_12_[9]  (.D(\sr_11_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[9]_net_1 ));
    DFN1E1C0 \sr_12_[11]  (.D(\sr_11_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[11]_net_1 ));
    DFN1E1C0 \sr_55_[9]  (.D(\sr_54_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[9]_net_1 ));
    DFN1E1C0 \sr_56_[8]  (.D(\sr_55_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[8]_net_1 ));
    DFN1E1C0 \sr_25_[6]  (.D(\sr_24_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[6]_net_1 ));
    DFN1E1C0 \sr_14_[3]  (.D(\sr_13_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[3]_net_1 ));
    DFN1E1C0 \sr_42_[0]  (.D(\sr_41_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[0]_net_1 ));
    DFN1E1C0 \sr_1_[7]  (.D(sr_new[7]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[7]));
    DFN1E1C0 \sr_2_[5]  (.D(sr_prev[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[5]_net_1 ));
    DFN1E1C0 \sr_14_[11]  (.D(\sr_13_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[11]_net_1 ));
    DFN1E1C0 \sr_37_[0]  (.D(\sr_36_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[0]_net_1 ));
    DFN1E1C0 \sr_58_[1]  (.D(\sr_57_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[1]_net_1 ));
    DFN1E1C0 \sr_11_[1]  (.D(\sr_10_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[1]_net_1 ));
    DFN1E1C0 \sr_62_[3]  (.D(\sr_61_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[3]_net_1 ));
    DFN1E1C0 \sr_45_[10]  (.D(\sr_44_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[10]_net_1 ));
    DFN1E1C0 \sr_16_[5]  (.D(\sr_15_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[5]_net_1 ));
    DFN1E1C0 \sr_43_[3]  (.D(\sr_42_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[3]_net_1 ));
    DFN1E1C0 \sr_61_[5]  (.D(\sr_60_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[5]_net_1 ));
    DFN1E1C0 \sr_54_[0]  (.D(\sr_53_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[0]_net_1 ));
    DFN1E1C0 \sr_16_[3]  (.D(\sr_15_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[3]_net_1 ));
    DFN1E1C0 \sr_4_[9]  (.D(\sr_3_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[9]_net_1 ));
    DFN1E1C0 \sr_40_[7]  (.D(\sr_39_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[7]_net_1 ));
    DFN1E1C0 \sr_50_[7]  (.D(\sr_49_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[7]_net_1 ));
    DFN1E1C0 \sr_31_[5]  (.D(\sr_30_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[5]_net_1 ));
    DFN1E1C0 \sr_50_[8]  (.D(\sr_49_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[8]_net_1 ));
    DFN1E1C0 \sr_49_[4]  (.D(\sr_48_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[4]_net_1 ));
    DFN1E1C0 \sr_31_[4]  (.D(\sr_30_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[4]_net_1 ));
    DFN1E1C0 \sr_0_[12]  (.D(cur_error[12]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable), .Q(sr_new[12]));
    DFN1E1C0 \sr_39_[3]  (.D(\sr_38_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[3]_net_1 ));
    DFN1E1C0 \sr_6_[7]  (.D(\sr_5_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[7]_net_1 ));
    DFN1E1C0 \sr_60_[7]  (.D(\sr_59_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[7]_net_1 ));
    DFN1E1C0 \sr_59_[6]  (.D(\sr_58_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[6]_net_1 ));
    DFN1E1C0 \sr_7_[3]  (.D(\sr_6_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[3]_net_1 ));
    DFN1E1C0 \sr_46_[10]  (.D(\sr_45_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[10]_net_1 ));
    DFN1E1C0 \sr_60_[8]  (.D(\sr_59_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[8]_net_1 ));
    DFN1E1C0 \sr_29_[4]  (.D(\sr_28_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[4]_net_1 ));
    DFN1E1C0 \sr_57_[11]  (.D(\sr_56_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[11]_net_1 ));
    DFN1E1C0 \sr_56_[0]  (.D(\sr_55_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[0]_net_1 ));
    DFN1E1C0 \sr_5_[7]  (.D(\sr_4_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[7]_net_1 ));
    DFN1E1C0 \sr_18_[7]  (.D(\sr_17_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[7]_net_1 ));
    DFN1E1C0 \sr_10_[5]  (.D(\sr_9_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[5]_net_1 ));
    DFN1E1C0 \sr_41_[12]  (.D(\sr_40_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[12]_net_1 ));
    DFN1E1C0 \sr_52_[10]  (.D(\sr_51_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[10]_net_1 ));
    DFN1E1C0 \sr_27_[11]  (.D(\sr_26_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[11]_net_1 ));
    DFN1E1C0 \sr_39_[12]  (.D(\sr_38_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[12]_net_1 ));
    DFN1E1C0 \sr_18_[6]  (.D(\sr_17_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_18_[6]_net_1 ));
    DFN1E1C0 \sr_22_[10]  (.D(\sr_21_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_22_[10]_net_1 ));
    DFN1E1C0 \sr_10_[3]  (.D(\sr_9_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[3]_net_1 ));
    DFN1E1C0 \sr_48_[5]  (.D(\sr_47_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[5]_net_1 ));
    DFN1E1C0 \sr_60_[0]  (.D(\sr_59_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[0]_net_1 ));
    DFN1E1C0 \sr_47_[4]  (.D(\sr_46_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[4]_net_1 ));
    DFN1E1C0 \sr_30_[12]  (.D(\sr_29_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[12]_net_1 ));
    DFN1E1C0 \sr_37_[3]  (.D(\sr_36_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[3]_net_1 ));
    DFN1E1C0 \sr_57_[6]  (.D(\sr_56_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[6]_net_1 ));
    DFN1E1C0 \sr_49_[6]  (.D(\sr_48_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[6]_net_1 ));
    DFN1E1C0 \sr_3_[3]  (.D(\sr_2_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[3]_net_1 ));
    DFN1E1C0 \sr_28_[9]  (.D(\sr_27_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[9]_net_1 ));
    DFN1E1C0 \sr_27_[4]  (.D(\sr_26_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[4]_net_1 ));
    DFN1E1C0 \sr_62_[12]  (.D(\sr_61_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[12]_net_1 ));
    DFN1E1C0 \sr_50_[0]  (.D(\sr_49_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[0]_net_1 ));
    DFN1E1C0 \sr_53_[9]  (.D(\sr_52_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[9]_net_1 ));
    DFN1E1C0 \sr_23_[6]  (.D(\sr_22_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[6]_net_1 ));
    DFN1E1C0 \sr_28_[1]  (.D(\sr_27_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[1]_net_1 ));
    DFN1E1C0 \sr_11_[4]  (.D(\sr_10_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[4]_net_1 ));
    DFN1E1C0 \sr_30_[10]  (.D(\sr_29_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[10]_net_1 ));
    DFN1E1C0 \sr_21_[8]  (.D(\sr_20_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[8]_net_1 ));
    DFN1E1C0 \sr_16_[12]  (.D(\sr_15_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[12]_net_1 ));
    DFN1E1C0 \sr_41_[10]  (.D(\sr_40_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[10]_net_1 ));
    DFN1E1C0 \sr_45_[1]  (.D(\sr_44_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[1]_net_1 ));
    DFN1E1C0 \sr_33_[10]  (.D(\sr_32_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[10]_net_1 ));
    DFN1E1C0 \sr_14_[12]  (.D(\sr_13_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[12]_net_1 ));
    DFN1E1C0 \sr_41_[11]  (.D(\sr_40_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[11]_net_1 ));
    DFN1E1C0 \sr_55_[12]  (.D(\sr_54_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[12]_net_1 ));
    DFN1E1C0 \sr_42_[7]  (.D(\sr_41_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[7]_net_1 ));
    DFN1E1C0 \sr_52_[7]  (.D(\sr_51_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[7]_net_1 ));
    DFN1E1C0 \sr_41_[2]  (.D(\sr_40_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[2]_net_1 ));
    DFN1E1C0 \sr_52_[8]  (.D(\sr_51_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[8]_net_1 ));
    DFN1E1C0 \sr_25_[12]  (.D(\sr_24_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[12]_net_1 ));
    DFN1E1C0 \sr_47_[6]  (.D(\sr_46_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[6]_net_1 ));
    DFN1E1C0 \sr_62_[7]  (.D(\sr_61_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[7]_net_1 ));
    DFN1E1C0 \sr_62_[8]  (.D(\sr_61_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[8]_net_1 ));
    DFN1E1C0 \sr_19_[1]  (.D(\sr_18_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[1]_net_1 ));
    DFN1E1C0 \sr_21_[0]  (.D(\sr_20_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[0]_net_1 ));
    DFN1E1C0 \sr_39_[10]  (.D(\sr_38_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[10]_net_1 ));
    DFN1E1C0 \sr_12_[5]  (.D(\sr_11_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[5]_net_1 ));
    DFN1E1C0 \sr_0_[10]  (.D(cur_error[10]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(int_enable), .Q(sr_new[10]));
    DFN1E1C0 \sr_12_[3]  (.D(\sr_11_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_12_[3]_net_1 ));
    DFN1E1C0 \sr_34_[1]  (.D(\sr_33_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[1]_net_1 ));
    DFN1E1C0 \sr_39_[5]  (.D(\sr_38_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[5]_net_1 ));
    DFN1E1C0 \sr_5_[11]  (.D(\sr_4_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[11]_net_1 ));
    DFN1E1C0 \sr_34_[2]  (.D(\sr_33_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[2]_net_1 ));
    DFN1E1C0 \sr_39_[4]  (.D(\sr_38_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[4]_net_1 ));
    DFN1E1C0 \sr_55_[2]  (.D(\sr_54_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[2]_net_1 ));
    DFN1E1C0 \sr_62_[0]  (.D(\sr_61_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[0]_net_1 ));
    DFN1E1C0 \sr_34_[7]  (.D(\sr_33_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[7]_net_1 ));
    DFN1E1C0 \sr_41_[8]  (.D(\sr_40_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_41_[8]_net_1 ));
    DFN1E1C0 \sr_52_[0]  (.D(\sr_51_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_52_[0]_net_1 ));
    DFN1E1C0 \sr_17_[1]  (.D(\sr_16_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[1]_net_1 ));
    DFN1E1C0 \sr_4_[0]  (.D(\sr_3_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[0]_net_1 ));
    DFN1E1C0 \sr_36_[1]  (.D(\sr_35_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[1]_net_1 ));
    DFN1E1C0 \sr_13_[12]  (.D(\sr_12_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[12]_net_1 ));
    DFN1E1C0 \sr_4_[6]  (.D(\sr_3_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[6]_net_1 ));
    DFN1E1C0 \sr_44_[9]  (.D(\sr_43_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[9]_net_1 ));
    DFN1E1C0 \sr_0_[3]  (.D(cur_error[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[3]));
    DFN1E1C0 \sr_36_[2]  (.D(\sr_35_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[2]_net_1 ));
    DFN1E1C0 \sr_51_[3]  (.D(\sr_50_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[3]_net_1 ));
    DFN1E1C0 \sr_36_[7]  (.D(\sr_35_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[7]_net_1 ));
    DFN1E1C0 \sr_21_[2]  (.D(\sr_20_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[2]_net_1 ));
    DFN1E1C0 \sr_37_[5]  (.D(\sr_36_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[5]_net_1 ));
    DFN1E1C0 \sr_55_[4]  (.D(\sr_54_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[4]_net_1 ));
    DFN1E1C0 \sr_21_[5]  (.D(\sr_20_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[5]_net_1 ));
    DFN1E1C0 \sr_43_[1]  (.D(\sr_42_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[1]_net_1 ));
    DFN1E1C0 \sr_11_[8]  (.D(\sr_10_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[8]_net_1 ));
    DFN1E1C0 \sr_37_[4]  (.D(\sr_36_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[4]_net_1 ));
    DFN1E1C0 \sr_62_[11]  (.D(\sr_61_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_62_[11]_net_1 ));
    DFN1E1C0 \sr_46_[9]  (.D(\sr_45_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[9]_net_1 ));
    DFN1E1C0 \sr_25_[7]  (.D(\sr_24_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[7]_net_1 ));
    DFN1E1C0 \sr_48_[3]  (.D(\sr_47_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[3]_net_1 ));
    DFN1E1C0 \sr_30_[1]  (.D(\sr_29_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[1]_net_1 ));
    DFN1E1C0 \sr_4_[1]  (.D(\sr_3_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[1]_net_1 ));
    DFN1E1C0 \sr_55_[10]  (.D(\sr_54_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[10]_net_1 ));
    DFN1E1C0 \sr_19_[4]  (.D(\sr_18_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[4]_net_1 ));
    DFN1E1C0 \sr_9_[7]  (.D(\sr_8_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[7]_net_1 ));
    DFN1E1C0 \sr_7_[4]  (.D(\sr_6_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[4]_net_1 ));
    DFN1E1C0 \sr_29_[8]  (.D(\sr_28_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[8]_net_1 ));
    DFN1E1C0 \sr_1_[3]  (.D(sr_new[3]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[3]));
    DFN1E1C0 \sr_34_[0]  (.D(\sr_33_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[0]_net_1 ));
    DFN1E1C0 \sr_30_[2]  (.D(\sr_29_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[2]_net_1 ));
    DFN1E1C0 \sr_25_[10]  (.D(\sr_24_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_25_[10]_net_1 ));
    DFN1E1C0 \sr_30_[7]  (.D(\sr_29_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[7]_net_1 ));
    DFN1E1C0 \sr_49_[2]  (.D(\sr_48_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[2]_net_1 ));
    DFN1E1C0 \sr_56_[10]  (.D(\sr_55_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[10]_net_1 ));
    DFN1E1C0 \sr_40_[9]  (.D(\sr_39_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[9]_net_1 ));
    DFN1E1C0 \sr_36_[0]  (.D(\sr_35_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[0]_net_1 ));
    DFN1E1C0 \sr_11_[2]  (.D(\sr_10_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[2]_net_1 ));
    DFN1E1C0 \sr_30_[11]  (.D(\sr_29_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[11]_net_1 ));
    DFN1E1C0 \sr_53_[2]  (.D(\sr_52_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[2]_net_1 ));
    DFN1E1C0 \sr_26_[10]  (.D(\sr_25_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[10]_net_1 ));
    DFN1E1C0 \sr_11_[0]  (.D(\sr_10_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[0]_net_1 ));
    DFN1E1C0 \sr_31_[8]  (.D(\sr_30_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[8]_net_1 ));
    DFN1E1C0 \sr_29_[0]  (.D(\sr_28_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[0]_net_1 ));
    DFN1E1C0 \sr_17_[4]  (.D(\sr_16_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[4]_net_1 ));
    DFN1E1C0 \sr_6_[3]  (.D(\sr_5_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[3]_net_1 ));
    DFN1E1C0 \sr_51_[12]  (.D(\sr_50_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[12]_net_1 ));
    DFN1E1C0 \sr_27_[8]  (.D(\sr_26_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[8]_net_1 ));
    DFN1E1C0 \sr_3_[4]  (.D(\sr_2_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[4]_net_1 ));
    DFN1E1C0 \sr_63_[2]  (.D(\sr_62_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[2]));
    DFN1E1C0 \sr_21_[12]  (.D(\sr_20_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[12]_net_1 ));
    DFN1E1C0 \sr_5_[3]  (.D(\sr_4_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_5_[3]_net_1 ));
    DFN1E1C0 \sr_15_[9]  (.D(\sr_14_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[9]_net_1 ));
    DFN1E1C0 \sr_51_[5]  (.D(\sr_50_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[5]_net_1 ));
    DFN1E1C0 \sr_47_[2]  (.D(\sr_46_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[2]_net_1 ));
    DFN1E1C0 \sr_47_[10]  (.D(\sr_46_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[10]_net_1 ));
    DFN1E1C0 \sr_45_[0]  (.D(\sr_44_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[0]_net_1 ));
    DFN1E1C0 \sr_58_[9]  (.D(\sr_57_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_58_[9]_net_1 ));
    DFN1E1C0 \sr_30_[0]  (.D(\sr_29_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[0]_net_1 ));
    DFN1E1C0 \sr_44_[4]  (.D(\sr_43_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[4]_net_1 ));
    DFN1E1C0 \sr_53_[4]  (.D(\sr_52_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_53_[4]_net_1 ));
    DFN1E1C0 \sr_34_[3]  (.D(\sr_33_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[3]_net_1 ));
    DFN1E1C0 \sr_54_[6]  (.D(\sr_53_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_54_[6]_net_1 ));
    DFN1E1C0 \sr_49_[8]  (.D(\sr_48_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[8]_net_1 ));
    DFN1E1C0 \sr_28_[6]  (.D(\sr_27_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_28_[6]_net_1 ));
    DFN1E1C0 \sr_21_[3]  (.D(\sr_20_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[3]_net_1 ));
    DFN1E1C0 \sr_31_[9]  (.D(\sr_30_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[9]_net_1 ));
    DFN1E1C0 \sr_8_[7]  (.D(\sr_7_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_8_[7]_net_1 ));
    DFN1E1C0 \sr_27_[0]  (.D(\sr_26_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[0]_net_1 ));
    DFN1E1C0 \sr_24_[4]  (.D(\sr_23_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_24_[4]_net_1 ));
    DFN1E1C0 \sr_63_[4]  (.D(\sr_62_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[4]));
    DFN1E1C0 \sr_32_[1]  (.D(\sr_31_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[1]_net_1 ));
    DFN1E1C0 \sr_19_[12]  (.D(\sr_18_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[12]_net_1 ));
    DFN1E1C0 \sr_23_[7]  (.D(\sr_22_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_23_[7]_net_1 ));
    DFN1E1C0 \sr_51_[10]  (.D(\sr_50_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[10]_net_1 ));
    DFN1E1C0 \sr_32_[2]  (.D(\sr_31_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[2]_net_1 ));
    DFN1E1C0 \sr_38_[12]  (.D(\sr_37_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[12]_net_1 ));
    DFN1E1C0 \sr_59_[3]  (.D(\sr_58_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[3]_net_1 ));
    DFN1E1C0 \sr_51_[11]  (.D(\sr_50_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[11]_net_1 ));
    DFN1E1C0 \sr_29_[2]  (.D(\sr_28_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[2]_net_1 ));
    DFN1E1C0 \sr_32_[7]  (.D(\sr_31_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[7]_net_1 ));
    DFN1E1C0 \sr_21_[10]  (.D(\sr_20_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[10]_net_1 ));
    DFN1E1C0 \sr_46_[4]  (.D(\sr_45_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[4]_net_1 ));
    DFN1E1C0 \sr_31_[6]  (.D(\sr_30_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_31_[6]_net_1 ));
    DFN1E1C0 \sr_36_[3]  (.D(\sr_35_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_36_[3]_net_1 ));
    DFN1E1C0 \sr_29_[5]  (.D(\sr_28_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[5]_net_1 ));
    DFN1E1C0 \sr_56_[6]  (.D(\sr_55_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_56_[6]_net_1 ));
    DFN1E1C0 \sr_21_[11]  (.D(\sr_20_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_21_[11]_net_1 ));
    DFN1E1C0 \sr_19_[8]  (.D(\sr_18_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[8]_net_1 ));
    DFN1E1C0 \sr_44_[10]  (.D(\sr_43_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[10]_net_1 ));
    DFN1E1C0 \sr_10_[12]  (.D(\sr_9_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[12]_net_1 ));
    DFN1E1C0 \sr_26_[4]  (.D(\sr_25_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_26_[4]_net_1 ));
    DFN1E1C0 \sr_47_[8]  (.D(\sr_46_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_47_[8]_net_1 ));
    DFN1E1C0 \sr_44_[6]  (.D(\sr_43_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_44_[6]_net_1 ));
    DFN1E1C0 \sr_42_[9]  (.D(\sr_41_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[9]_net_1 ));
    DFN1E1C0 \sr_63_[9]  (.D(\sr_62_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[9]));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \sr_10_[10]  (.D(\sr_9_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_10_[10]_net_1 ));
    DFN1E1C0 \sr_2_[10]  (.D(sr_prev[10]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[10]_net_1 ));
    DFN1E1C0 \sr_13_[10]  (.D(\sr_12_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[10]_net_1 ));
    DFN1E1C0 \sr_57_[3]  (.D(\sr_56_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_57_[3]_net_1 ));
    DFN1E1C0 \sr_27_[2]  (.D(\sr_26_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[2]_net_1 ));
    DFN1E1C0 \sr_40_[4]  (.D(\sr_39_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[4]_net_1 ));
    DFN1E1C0 \sr_30_[3]  (.D(\sr_29_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_30_[3]_net_1 ));
    DFN1E1C0 \sr_50_[6]  (.D(\sr_49_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_50_[6]_net_1 ));
    DFN1E1C0 \sr_27_[5]  (.D(\sr_26_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_27_[5]_net_1 ));
    DFN1E1C0 \sr_46_[6]  (.D(\sr_45_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[6]_net_1 ));
    DFN1E1C0 \sr_38_[11]  (.D(\sr_37_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_38_[11]_net_1 ));
    DFN1E1C0 \sr_17_[8]  (.D(\sr_16_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[8]_net_1 ));
    DFN1E1C0 \sr_20_[4]  (.D(\sr_19_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_20_[4]_net_1 ));
    DFN1E1C0 \sr_0_[4]  (.D(cur_error[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(sr_new[4]));
    DFN1E1C0 \sr_49_[11]  (.D(\sr_48_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_49_[11]_net_1 ));
    DFN1E1C0 \sr_13_[9]  (.D(\sr_12_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_13_[9]_net_1 ));
    DFN1E1C0 \sr_60_[6]  (.D(\sr_59_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_60_[6]_net_1 ));
    DFN1E1C0 \sr_2_[7]  (.D(sr_prev[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(int_enable), .Q(\sr_2_[7]_net_1 ));
    DFN1E1C0 \sr_51_[1]  (.D(\sr_50_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_51_[1]_net_1 ));
    DFN1E1C0 \sr_32_[0]  (.D(\sr_31_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_32_[0]_net_1 ));
    DFN1E1C0 \sr_7_[2]  (.D(\sr_6_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[2]_net_1 ));
    DFN1E1C0 \sr_4_[11]  (.D(\sr_3_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[11]_net_1 ));
    DFN1E1C0 \sr_19_[2]  (.D(\sr_18_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[2]_net_1 ));
    DFN1E1C0 \sr_7_[8]  (.D(\sr_6_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_7_[8]_net_1 ));
    DFN1E1C0 \sr_4_[5]  (.D(\sr_3_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_4_[5]_net_1 ));
    DFN1E1C0 \sr_43_[0]  (.D(\sr_42_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_43_[0]_net_1 ));
    DFN1E1C0 \sr_19_[0]  (.D(\sr_18_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[0]_net_1 ));
    DFN1E1C0 \sr_9_[10]  (.D(\sr_8_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_9_[10]_net_1 ));
    DFN1E1C0 \sr_39_[8]  (.D(\sr_38_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[8]_net_1 ));
    DFN1E1C0 \sr_61_[1]  (.D(\sr_60_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_61_[1]_net_1 ));
    DFN1E1C0 \sr_19_[10]  (.D(\sr_18_[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_19_[10]_net_1 ));
    DFN1E1C0 \sr_14_[1]  (.D(\sr_13_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_14_[1]_net_1 ));
    DFN1E1C0 \sr_63_[3]  (.D(\sr_62_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[3]));
    DFN1E1C0 \sr_45_[7]  (.D(\sr_44_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_45_[7]_net_1 ));
    DFN1E1C0 \sr_59_[5]  (.D(\sr_58_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_59_[5]_net_1 ));
    DFN1E1C0 \sr_55_[7]  (.D(\sr_54_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[7]_net_1 ));
    DFN1E1C0 \sr_63_[12]  (.D(\sr_62_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(sr_old[12]));
    DFN1E1C0 \sr_48_[1]  (.D(\sr_47_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_48_[1]_net_1 ));
    DFN1E1C0 \sr_42_[12]  (.D(\sr_41_[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_42_[12]_net_1 ));
    DFN1E1C0 \sr_40_[6]  (.D(\sr_39_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_40_[6]_net_1 ));
    DFN1E1C0 \sr_55_[8]  (.D(\sr_54_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_55_[8]_net_1 ));
    DFN1E1C0 \sr_1_[4]  (.D(sr_new[4]), .CLK(clk_c), .CLR(n_rst_c), .E(
        int_enable), .Q(sr_prev[4]));
    DFN1E1C0 \sr_34_[5]  (.D(\sr_33_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[5]_net_1 ));
    DFN1E1C0 \sr_6_[11]  (.D(\sr_5_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_6_[11]_net_1 ));
    DFN1E1C0 \sr_11_[7]  (.D(\sr_10_[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[7]_net_1 ));
    DFN1E1C0 \sr_34_[4]  (.D(\sr_33_[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_34_[4]_net_1 ));
    DFN1E1C0 \sr_16_[1]  (.D(\sr_15_[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_16_[1]_net_1 ));
    DFN1E1C0 \sr_29_[3]  (.D(\sr_28_[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_29_[3]_net_1 ));
    DFN1E1C0 \sr_17_[2]  (.D(\sr_16_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[2]_net_1 ));
    DFN1E1C0 \sr_39_[9]  (.D(\sr_38_[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_39_[9]_net_1 ));
    DFN1E1C0 \sr_3_[2]  (.D(\sr_2_[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[2]_net_1 ));
    DFN1E1C0 \sr_46_[11]  (.D(\sr_45_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_46_[11]_net_1 ));
    DFN1E1C0 \sr_3_[8]  (.D(\sr_2_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_3_[8]_net_1 ));
    DFN1E1C0 \sr_33_[11]  (.D(\sr_32_[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_33_[11]_net_1 ));
    DFN1E1C0 \sr_17_[0]  (.D(\sr_16_[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_17_[0]_net_1 ));
    DFN1E1C0 \sr_37_[8]  (.D(\sr_36_[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_37_[8]_net_1 ));
    DFN1E1C0 \sr_15_[5]  (.D(\sr_14_[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_15_[5]_net_1 ));
    DFN1E1C0 \sr_11_[6]  (.D(\sr_10_[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(int_enable), .Q(\sr_11_[6]_net_1 ));
    
endmodule


module controller_Z1_4_3(
       pwm_chg,
       N_46_1_0,
       N_46_1,
       sig_prev_0,
       sig_old_i_0_0,
       pwm_rdy,
       sig_old_i_0,
       sig_prev,
       sum_rdy,
       deriv_enable,
       calc_avg,
       calc_int,
       pwm_enable,
       sum_enable,
       calc_error,
       avg_enable,
       int_enable,
       pwm_chg_0,
       avg_enable_0,
       n_rst_c,
       clk_c,
       avg_enable_1
    );
output pwm_chg;
input  N_46_1_0;
input  N_46_1;
input  sig_prev_0;
input  sig_old_i_0_0;
input  pwm_rdy;
input  sig_old_i_0;
input  sig_prev;
input  sum_rdy;
output deriv_enable;
output calc_avg;
output calc_int;
output pwm_enable;
output sum_enable;
output calc_error;
output avg_enable;
output int_enable;
output pwm_chg_0;
output avg_enable_0;
input  n_rst_c;
input  clk_c;
output avg_enable_1;

    wire \state_RNIIJEQ2[0]_net_1 , N_12, \state_2[5] , N_94, 
        \count[13]_net_1 , count_c12, count_31_0, count_n14, 
        count_n14_tz, N_62, \count[14]_net_1 , count_n13, count_n12, 
        count_c11, \count[12]_net_1 , count_n11, count_c10, 
        \count[11]_net_1 , count_n15, \count[15]_net_1 , count_c9, 
        \count[10]_net_1 , count_c8, \count[9]_net_1 , count_c7, 
        \count[8]_net_1 , count_c6, \count[7]_net_1 , count_c5, 
        \count[6]_net_1 , count_c4, \count[5]_net_1 , count_c3, 
        \count[4]_net_1 , count_c2, \count[3]_net_1 , count_c1, 
        \count[0]_net_1 , \count[1]_net_1 , \count[2]_net_1 , 
        \state_ns_0_a2_9[0] , \state[10]_net_1 , N_33, 
        \state_ns_0_a2_8[0] , \state_ns_0_a2_6[0] , 
        \state_ns_0_a2_5[0] , \state_ns_0_a2_2[0] , N_270, N_272, 
        \state_ns_0_a2_1[0] , \state_ns_0_a2_0[0] , \state[7]_net_1 , 
        next_state_0_sqmuxa_1_1_a2_0_a2_0, \state_ns_i_0_0[2] , 
        un1_countlto15_13, un1_countlto15_5, un1_countlto15_4, 
        un1_countlto15_11, un1_countlto15_12, un1_countlto15_1, 
        un1_countlto15_0, un1_countlto15_9, un1_countlto15_7, 
        un1_countlto15_3, N_274, N_23, N_273, \state[0]_net_1 , N_26, 
        next_state15_li, \state_RNIEUBQ[4]_net_1 , \state_RNO_2[5] , 
        N_24, count_n10, count_n9, count_n2, count_n3, count_n4, 
        count_n5, count_n6, count_n7, count_n8, \state[4]_net_1 , 
        \state[12]_net_1 , count_n1, N_267, \state_ns[12] , counte, 
        \state_RNO_3[8] , \state_ns[0] , \state_ns[1] , 
        \avg_count[1]_net_1 , \avg_count[0]_net_1 , \state_ns[7] , 
        \state_ns[10] , \state_ns[4] , \DWACT_ADD_CI_0_partial_sum[0] , 
        I_10_3, \DWACT_ADD_CI_0_TMP[0] , GND, VCC;
    
    DFN1E1C0 \count[5]  (.D(count_n5), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[5]_net_1 ));
    OA1A \state_RNO_0[0]  (.A(\state[10]_net_1 ), .B(N_33), .C(
        \state_ns_0_a2_8[0] ), .Y(\state_ns_0_a2_9[0] ));
    NOR3C \count_RNIS1S32[3]  (.A(un1_countlto15_5), .B(
        un1_countlto15_4), .C(un1_countlto15_11), .Y(un1_countlto15_13)
        );
    NOR2B \count_RNI94DA1[4]  (.A(count_c3), .B(\count[4]_net_1 ), .Y(
        count_c4));
    DFN1E1C0 \count[1]  (.D(count_n1), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[1]_net_1 ));
    DFN1E1C0 \count[10]  (.D(count_n10), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[10]_net_1 ));
    DFN1E1C0 \count[0]  (.D(N_267), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[0]_net_1 ));
    NOR2 \state_RNO_9[0]  (.A(calc_avg), .B(deriv_enable), .Y(
        \state_ns_0_a2_0[0] ));
    DFN1C0 \state[13]  (.D(N_12), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_chg));
    DFN1E1C0 \count[14]  (.D(count_n14), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[14]_net_1 ));
    DFN1C0 \state[7]  (.D(\state_ns[7] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[7]_net_1 ));
    AX1C \count_RNO_0[14]  (.A(\count[13]_net_1 ), .B(count_c12), .C(
        \count[14]_net_1 ), .Y(count_n14_tz));
    NOR3 \state_RNIIJEQ2[0]  (.A(N_274), .B(\state_ns_i_0_0[2] ), .C(
        N_23), .Y(\state_RNIIJEQ2[0]_net_1 ));
    NOR2B \count_RNIKPR32[7]  (.A(count_c6), .B(\count[7]_net_1 ), .Y(
        count_c7));
    NOR2B \count_RNIFNLS2[10]  (.A(count_c9), .B(\count[10]_net_1 ), 
        .Y(count_c10));
    NOR2B \count_RNI7OUG[1]  (.A(\count[0]_net_1 ), .B(
        \count[1]_net_1 ), .Y(count_c1));
    DFN1C0 \state[5]  (.D(\state_RNO_2[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state_2[5] ));
    XA1B \count_RNO[7]  (.A(count_c6), .B(\count[7]_net_1 ), .C(N_62), 
        .Y(count_n7));
    AX1 \count_RNO[15]  (.A(N_62), .B(\count[15]_net_1 ), .C(N_94), .Y(
        count_n15));
    DFN1C0 \state[4]  (.D(\state_ns[4] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[4]_net_1 ));
    XA1B \count_RNO[2]  (.A(count_c1), .B(\count[2]_net_1 ), .C(N_62), 
        .Y(count_n2));
    AO1A \state_RNO[7]  (.A(N_46_1), .B(\state[7]_net_1 ), .C(calc_int)
        , .Y(\state_ns[7] ));
    DFN1C0 \state_1[2]  (.D(\state_RNIIJEQ2[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable_1));
    NOR2B \count_RNIKDG43[11]  (.A(count_c10), .B(\count[11]_net_1 ), 
        .Y(count_c11));
    NOR2A \state_RNO_0[5]  (.A(N_272), .B(\state[10]_net_1 ), .Y(N_24));
    DFN1C0 \state_0[2]  (.D(\state_RNIIJEQ2[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable_0));
    XA1B \count_RNO[9]  (.A(count_c8), .B(\count[9]_net_1 ), .C(N_62), 
        .Y(count_n9));
    OR2B \state_RNID8KH[4]  (.A(\state[4]_net_1 ), .B(
        \state[12]_net_1 ), .Y(N_273));
    DFN1C0 \state[6]  (.D(int_enable), .CLK(clk_c), .CLR(n_rst_c), .Q(
        calc_int));
    NOR2B \count_RNIB2RK2[9]  (.A(count_c8), .B(\count[9]_net_1 ), .Y(
        count_c9));
    NOR2 \state_RNO_6[0]  (.A(sum_enable), .B(\state[7]_net_1 ), .Y(
        \state_ns_0_a2_2[0] ));
    DFN1C0 \state[2]  (.D(\state_RNIIJEQ2[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(avg_enable));
    VCC VCC_i (.Y(VCC));
    XOR2 un1_avg_count_1_I_10 (.A(\avg_count[1]_net_1 ), .B(
        \DWACT_ADD_CI_0_TMP[0] ), .Y(I_10_3));
    XA1B \count_RNO[4]  (.A(count_c3), .B(\count[4]_net_1 ), .C(N_62), 
        .Y(count_n4));
    DFN1C0 \state[3]  (.D(avg_enable), .CLK(clk_c), .CLR(n_rst_c), .Q(
        calc_avg));
    DFN1E1C0 \count[8]  (.D(count_n8), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[8]_net_1 ));
    NOR2B \state_RNIPGSS[12]  (.A(pwm_rdy), .B(\state[12]_net_1 ), .Y(
        N_12));
    NOR2 \count_RNIFHLF[14]  (.A(\count[14]_net_1 ), .B(
        \count[13]_net_1 ), .Y(un1_countlto15_1));
    XA1B \count_RNO[10]  (.A(count_c9), .B(\count[10]_net_1 ), .C(N_62)
        , .Y(count_n10));
    NOR2B \state_RNO[8]  (.A(\state[7]_net_1 ), .B(N_46_1), .Y(
        \state_RNO_3[8] ));
    NOR3B \state_RNO_1[0]  (.A(next_state15_li), .B(
        \state_RNIEUBQ[4]_net_1 ), .C(\state[10]_net_1 ), .Y(N_26));
    DFN1E1C0 \count[15]  (.D(count_n15), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[15]_net_1 ));
    XA1B \count_RNO[3]  (.A(count_c2), .B(\count[3]_net_1 ), .C(N_62), 
        .Y(count_n3));
    NOR2B \count_RNI1LSI1[5]  (.A(count_c4), .B(\count[5]_net_1 ), .Y(
        count_c5));
    DFN1E1C0 \count[11]  (.D(count_n11), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[11]_net_1 ));
    NOR2B \state_RNIEUBQ[4]  (.A(\state[4]_net_1 ), .B(N_46_1_0), .Y(
        \state_RNIEUBQ[4]_net_1 ));
    DFN1C0 \state_0[13]  (.D(N_12), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_chg_0));
    XA1B \count_RNO[8]  (.A(count_c7), .B(\count[8]_net_1 ), .C(N_62), 
        .Y(count_n8));
    OR2B \avg_count_RNI1UVM[1]  (.A(\avg_count[1]_net_1 ), .B(
        \avg_count[0]_net_1 ), .Y(next_state15_li));
    AO1A \state_RNO[10]  (.A(sum_rdy), .B(\state[10]_net_1 ), .C(
        sum_enable), .Y(\state_ns[10] ));
    NOR2B \count_RNIIKT11[3]  (.A(count_c2), .B(\count[3]_net_1 ), .Y(
        count_c3));
    DFN1E1C0 \count[13]  (.D(count_n13), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[13]_net_1 ));
    XA1B \count_RNO[5]  (.A(count_c4), .B(\count[5]_net_1 ), .C(N_62), 
        .Y(count_n5));
    XA1B \count_RNO[1]  (.A(\count[1]_net_1 ), .B(\count[0]_net_1 ), 
        .C(N_62), .Y(count_n1));
    XA1B \count_RNO[11]  (.A(count_c10), .B(\count[11]_net_1 ), .C(
        N_62), .Y(count_n11));
    NOR2 \count_RNIL6VG[7]  (.A(\count[7]_net_1 ), .B(\count[8]_net_1 )
        , .Y(un1_countlto15_4));
    NOR3A \count_RNIMOT11[3]  (.A(un1_countlto15_7), .B(
        \count[4]_net_1 ), .C(\count[3]_net_1 ), .Y(un1_countlto15_11));
    NOR3B \state_RNO_4[0]  (.A(\state_ns_0_a2_2[0] ), .B(N_270), .C(
        N_272), .Y(\state_ns_0_a2_6[0] ));
    DFN1C0 \state[11]  (.D(N_62), .CLK(clk_c), .CLR(n_rst_c), .Q(
        pwm_enable));
    DFN1E1C0 \count[2]  (.D(count_n2), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[2]_net_1 ));
    NOR2 \count_RNI0AAG[10]  (.A(\count[10]_net_1 ), .B(
        \count[9]_net_1 ), .Y(un1_countlto15_3));
    DFN1P0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .PRE(n_rst_c), 
        .Q(\state[0]_net_1 ));
    DFN1C0 \state[12]  (.D(\state_ns[12] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[12]_net_1 ));
    NOR2A \count_RNO_1[15]  (.A(\count[14]_net_1 ), .B(N_62), .Y(
        count_31_0));
    NOR2B \count_RNIS5EP[2]  (.A(count_c1), .B(\count[2]_net_1 ), .Y(
        count_c2));
    GND GND_i (.Y(GND));
    NOR3A \count_RNIBNVV[11]  (.A(un1_countlto15_3), .B(
        \count[11]_net_1 ), .C(\count[12]_net_1 ), .Y(un1_countlto15_9)
        );
    DFN1E1C0 \count[9]  (.D(count_n9), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[9]_net_1 ));
    XA1B \count_RNO[6]  (.A(count_c5), .B(\count[6]_net_1 ), .C(N_62), 
        .Y(count_n6));
    XA1B \count_RNO[12]  (.A(count_c11), .B(\count[12]_net_1 ), .C(
        N_62), .Y(count_n12));
    NOR2 \count_RNO[0]  (.A(\count[0]_net_1 ), .B(N_62), .Y(N_267));
    AND2 un1_avg_count_1_I_1 (.A(\avg_count[0]_net_1 ), .B(
        \state_RNIEUBQ[4]_net_1 ), .Y(\DWACT_ADD_CI_0_TMP[0] ));
    XOR2 un1_avg_count_1_I_8 (.A(\avg_count[0]_net_1 ), .B(
        \state_RNIEUBQ[4]_net_1 ), .Y(\DWACT_ADD_CI_0_partial_sum[0] ));
    NOR3B \state_RNO_5[0]  (.A(\state_ns_0_a2_1[0] ), .B(
        \state_ns_0_a2_0[0] ), .C(calc_error), .Y(\state_ns_0_a2_5[0] )
        );
    NOR3C \state_RNO_2[0]  (.A(un1_countlto15_12), .B(
        un1_countlto15_13), .C(sum_rdy), .Y(N_33));
    NOR3A \state_RNIKA831[0]  (.A(N_273), .B(\state[10]_net_1 ), .C(
        \state[0]_net_1 ), .Y(N_274));
    AO1A \state_RNO[4]  (.A(N_46_1_0), .B(\state[4]_net_1 ), .C(
        calc_avg), .Y(\state_ns[4] ));
    CLKINT \state_RNIG5Q3[5]  (.A(\state_2[5] ), .Y(int_enable));
    NOR2 \count_RNIH2VG[5]  (.A(\count[5]_net_1 ), .B(\count[6]_net_1 )
        , .Y(un1_countlto15_5));
    NOR2B \count_RNIFDBC2[8]  (.A(count_c7), .B(\count[8]_net_1 ), .Y(
        count_c8));
    DFN1E1C0 \count[6]  (.D(count_n6), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[6]_net_1 ));
    AO1A \state_RNO[12]  (.A(pwm_rdy), .B(\state[12]_net_1 ), .C(
        pwm_enable), .Y(\state_ns[12] ));
    DFN1C0 \state[10]  (.D(\state_ns[10] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\state[10]_net_1 ));
    OR2 \state_RNID8KH_0[4]  (.A(\state[4]_net_1 ), .B(
        \state[12]_net_1 ), .Y(N_272));
    DFN1E1C0 \count[3]  (.D(count_n3), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[3]_net_1 ));
    DFN1C0 \state[1]  (.D(\state_ns[1] ), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(calc_error));
    NOR2 \state_RNO_8[0]  (.A(pwm_enable), .B(calc_int), .Y(
        \state_ns_0_a2_1[0] ));
    DFN1C0 \state[8]  (.D(\state_RNO_3[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(deriv_enable));
    NOR2B \count_RNIQ6CR1[6]  (.A(count_c5), .B(\count[6]_net_1 ), .Y(
        count_c6));
    NOR3C \count_RNIMEVV1[11]  (.A(un1_countlto15_1), .B(
        un1_countlto15_0), .C(un1_countlto15_9), .Y(un1_countlto15_12));
    NOR3A \state_RNO[5]  (.A(calc_error), .B(\state[7]_net_1 ), .C(
        N_24), .Y(\state_RNO_2[5] ));
    NOR2A \count_RNO[14]  (.A(count_n14_tz), .B(N_62), .Y(count_n14));
    NOR2B \state_RNIOHKM[10]  (.A(\state[10]_net_1 ), .B(sum_rdy), .Y(
        next_state_0_sqmuxa_1_1_a2_0_a2_0));
    XA1B \count_RNO[13]  (.A(count_c12), .B(\count[13]_net_1 ), .C(
        N_62), .Y(count_n13));
    DFN1C0 \state[9]  (.D(deriv_enable), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(sum_enable));
    NOR2 \count_RNI9QUG[1]  (.A(\count[1]_net_1 ), .B(\count[2]_net_1 )
        , .Y(un1_countlto15_7));
    NOR2 \state_RNIO8EL[0]  (.A(\state[0]_net_1 ), .B(N_272), .Y(N_23));
    DFN1C0 \avg_count[0]  (.D(\DWACT_ADD_CI_0_partial_sum[0] ), .CLK(
        clk_c), .CLR(n_rst_c), .Q(\avg_count[0]_net_1 ));
    OR3C \state_RNO_7[0]  (.A(sig_prev), .B(sig_old_i_0), .C(
        \state[0]_net_1 ), .Y(N_270));
    AO1A \state_RNO[0]  (.A(int_enable), .B(\state_ns_0_a2_9[0] ), .C(
        N_26), .Y(\state_ns[0] ));
    OR3B \state_RNI60O11[7]  (.A(sig_prev), .B(sig_old_i_0), .C(
        \state[7]_net_1 ), .Y(\state_ns_i_0_0[2] ));
    NOR2 \count_RNIS5AG[15]  (.A(\count[15]_net_1 ), .B(
        \count[0]_net_1 ), .Y(un1_countlto15_0));
    DFN1C0 \avg_count[1]  (.D(I_10_3), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \avg_count[1]_net_1 ));
    AOI1B \state_RNIA2GQ4[10]  (.A(un1_countlto15_13), .B(
        un1_countlto15_12), .C(next_state_0_sqmuxa_1_1_a2_0_a2_0), .Y(
        N_62));
    NOR3C \count_RNO_0[15]  (.A(\count[13]_net_1 ), .B(count_c12), .C(
        count_31_0), .Y(N_94));
    NOR2B \count_RNIQ4BC3[12]  (.A(count_c11), .B(\count[12]_net_1 ), 
        .Y(count_c12));
    NOR3B \state_RNO_3[0]  (.A(\state_ns_0_a2_6[0] ), .B(
        \state_ns_0_a2_5[0] ), .C(avg_enable), .Y(\state_ns_0_a2_8[0] )
        );
    AO1 \state_RNIAD6J5[10]  (.A(sig_old_i_0_0), .B(sig_prev_0), .C(
        N_62), .Y(counte));
    DFN1E1C0 \count[4]  (.D(count_n4), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[4]_net_1 ));
    DFN1E1C0 \count[12]  (.D(count_n12), .CLK(clk_c), .CLR(n_rst_c), 
        .E(counte), .Q(\count[12]_net_1 ));
    NOR2A \state_RNO[1]  (.A(\state_RNIEUBQ[4]_net_1 ), .B(
        next_state15_li), .Y(\state_ns[1] ));
    DFN1E1C0 \count[7]  (.D(count_n7), .CLK(clk_c), .CLR(n_rst_c), .E(
        counte), .Q(\count[7]_net_1 ));
    
endmodule


module sig_gen_8(
       primary_15_c,
       n_rst_c,
       clk_c,
       sig_old_i_0,
       sig_prev
    );
input  primary_15_c;
input  n_rst_c;
input  clk_c;
output sig_old_i_0;
output sig_prev;

    wire sig_prev_i, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(clk_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev_inst_1 (.D(primary_15_c), .CLK(clk_c), .CLR(
        n_rst_c), .Q(sig_prev));
    INV sig_old_RNO (.A(sig_prev), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module pid_sum_13s_4_3(
       integral_i,
       integral,
       derivative_0,
       sr_new,
       sr_new_0_0,
       integral_0_0,
       integral_1_0,
       sum_39,
       sum_14,
       sum_20,
       sum_19,
       sum_22,
       sum_13,
       sum_17,
       sum_18,
       sum_23,
       sum_21,
       sum_16,
       sum_15,
       sum_12,
       sum_11,
       sum_6,
       sum_9,
       sum_10,
       sum_5,
       sum_8,
       sum_7,
       sum_4,
       sum_2_d0,
       sum_1_d0,
       sum_0_d0,
       sum_3,
       sum_0_0,
       sum_1_0,
       sum_2_0,
       sum_enable,
       sum_rdy,
       n_rst_c,
       clk_c
    );
input  [25:24] integral_i;
input  [25:6] integral;
input  derivative_0;
input  [12:0] sr_new;
input  sr_new_0_0;
input  integral_0_0;
input  integral_1_0;
output sum_39;
output sum_14;
output sum_20;
output sum_19;
output sum_22;
output sum_13;
output sum_17;
output sum_18;
output sum_23;
output sum_21;
output sum_16;
output sum_15;
output sum_12;
output sum_11;
output sum_6;
output sum_9;
output sum_10;
output sum_5;
output sum_8;
output sum_7;
output sum_4;
output sum_2_d0;
output sum_1_d0;
output sum_0_d0;
output sum_3;
output sum_0_0;
output sum_1_0;
output sum_2_0;
input  sum_enable;
output sum_rdy;
input  n_rst_c;
input  clk_c;

    wire \next_sum[39] , N_416, \state_0[1]_net_1 , 
        \state_RNIGPKC[0]_net_1 , \state_2[2]_net_1 , 
        \state_1[2]_net_1 , \state_0[2]_net_1 , \state_0[3]_net_1 , 
        \state[6]_net_1 , N_416_0, \un1_next_sum_1_iv_0[26] , 
        next_sum_1_sqmuxa_2, next_sum_1_sqmuxa_1, next_sum_1_sqmuxa, 
        N_12, N_10, \DWACT_FINC_E[0] , N_5, \DWACT_FINC_E[4] , N_2, 
        \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , N_25, N_23, 
        \DWACT_FINC_E_0[0] , N_18, \DWACT_FINC_E_0[4] , N_15, 
        \DWACT_FINC_E_0[7] , \DWACT_FINC_E_0[6] , \un1_next_sum[21] , 
        N_228_1, \un1_next_sum_iv_0[21]_net_1 , \un1_next_sum[19] , 
        \un1_next_sum_iv_0[19]_net_1 , N586, \un1_next_sum_1_iv[26] , 
        \sumreg[38]_net_1 , \ireg_m[19] , \ireg[19]_net_1 , 
        \ireg_m[21] , \ireg[21]_net_1 , ADD_40x40_fast_I195_Y_1, N595, 
        ADD_40x40_fast_I195_Y_0, N583, \un3_next_sum_m[19] , 
        \un3_next_sum_m[21] , ADD_40x40_fast_I448_Y_0, 
        \sumreg[30]_net_1 , ADD_40x40_fast_I447_Y_0, 
        \sumreg[29]_net_1 , ADD_40x40_fast_I456_Y_0, 
        ADD_40x40_fast_I449_Y_0, \sumreg[31]_net_1 , 
        ADD_40x40_fast_I453_Y_0, \sumreg[35]_net_1 , 
        ADD_40x40_fast_I454_Y_0, \sumreg[36]_net_1 , 
        ADD_40x40_fast_I455_Y_0, \sumreg[37]_net_1 , 
        ADD_40x40_fast_I452_Y_0, \sumreg[34]_net_1 , 
        ADD_40x40_fast_I451_Y_0, \sumreg[33]_net_1 , 
        ADD_40x40_fast_I347_Y_0, N787, N772, N771, 
        ADD_40x40_fast_I457_Y_0, ADD_40x40_fast_I446_Y_0, 
        \sumreg[28]_net_1 , ADD_40x40_fast_I450_Y_0, 
        \sumreg[32]_net_1 , ADD_40x40_fast_I379_Y_4, N840, N871, 
        ADD_40x40_fast_I379_Y_3, N756, ADD_40x40_fast_I379_Y_2, N596, 
        ADD_40x40_fast_I379_Y_0, N681, ADD_40x40_fast_I346_Y_0, N785, 
        N770, N769, ADD_40x40_fast_I381_Y_2, N760, N775, 
        ADD_40x40_fast_I381_Y_1, N600, N685, ADD_40x40_fast_I382_Y_1, 
        N762, N777, ADD_40x40_fast_I382_Y_0, N598, N602, N687, 
        ADD_40x40_fast_I445_Y_0, \sumreg[27]_net_1 , 
        ADD_40x40_fast_I432_Y_0, \un1_next_sum[14] , 
        ADD_40x40_fast_I380_Y_2, N758, N773, ADD_40x40_fast_I380_Y_1, 
        N594, N683, ADD_40x40_fast_I347_un1_Y_0, N788, 
        ADD_40x40_fast_I438_Y_0, \un1_next_sum_iv_0[20] , 
        ADD_40x40_fast_I437_Y_0, ADD_40x40_fast_I384_Y_2, 
        ADD_40x40_fast_I384_Y_0, I278_un1_Y, I384_un1_Y, N691, N684, 
        ADD_40x40_fast_I383_Y_1, N764, N779, ADD_40x40_fast_I383_Y_0, 
        N608, N612, ADD_40x40_fast_I444_Y_0, \sumreg[26]_net_1 , 
        ADD_40x40_fast_I443_Y_0, \sumreg[25]_net_1 , 
        \un1_next_sum_0_iv[25] , ADD_40x40_fast_I440_Y_0, 
        \un1_next_sum[22] , ADD_40x40_fast_I378_Y_3, N754, 
        ADD_40x40_fast_I378_Y_2, ADD_40x40_fast_I378_Y_1, 
        ADD_40x40_fast_I378_Y_0, ADD_40x40_fast_I349_Y_0, N791, N776, 
        ADD_40x40_fast_I385_Y_1, N768, N783, ADD_40x40_fast_I385_Y_0, 
        I208_un1_Y, ADD_40x40_fast_I431_Y_0, \un1_next_sum[13] , 
        ADD_40x40_fast_I442_Y_0, \sumreg[24]_net_1 , 
        \un1_next_sum[24] , ADD_40x40_fast_I435_Y_0, 
        \un1_next_sum[17] , ADD_40x40_fast_I436_Y_0, 
        \un1_next_sum[18] , ADD_40x40_fast_I441_Y_0, 
        \un1_next_sum_iv_0[23] , ADD_40x40_fast_I439_Y_0, 
        ADD_40x40_fast_I434_Y_0, \un1_next_sum_iv_1[16] , 
        \un1_next_sum_iv_2[16] , ADD_40x40_fast_I433_Y_0, 
        \un1_next_sum[15] , ADD_40x40_fast_I346_un1_Y_0, N786, 
        ADD_40x40_fast_I430_Y_0, \un1_next_sum[12] , 
        ADD_40x40_fast_I349_un1_Y_0, N792, ADD_40x40_fast_I379_un1_Y_0, 
        N872, ADD_40x40_fast_I429_Y_0, \un1_next_sum_iv_1[11] , 
        \un1_next_sum_iv_2[11] , ADD_40x40_fast_I424_Y_0, 
        \un1_next_sum[6] , ADD_40x40_fast_I427_Y_0, 
        \un1_next_sum_iv_1[9] , \un1_next_sum_iv_2[9] , 
        ADD_40x40_fast_I428_Y_0, \un1_next_sum[10] , 
        ADD_40x40_fast_I352_un1_Y_0, N798, N782, 
        ADD_40x40_fast_I351_un1_Y_0, N706, N698, N796, 
        ADD_40x40_fast_I423_Y_0, \un1_next_sum_iv_0[5] , 
        ADD_40x40_fast_I426_Y_0, \un1_next_sum[8] , 
        ADD_40x40_fast_I353_un1_Y_0, N800, N784, 
        ADD_40x40_fast_I425_Y_0, \un1_next_sum[7] , 
        ADD_40x40_fast_I422_Y_0, \un1_next_sum[4] , 
        ADD_40x40_fast_I420_Y_0, \un1_next_sum[0] , 
        ADD_40x40_fast_I419_Y_0, ADD_40x40_fast_I257_Y_1, N475, N472, 
        N661, ADD_40x40_fast_I199_Y_0, N599, ADD_40x40_fast_I197_Y_0, 
        ADD_22x22_fast_I176_Y_0, \i_adj[18]_net_1 , \i_adj[16]_net_1 , 
        ADD_22x22_fast_I126_Y_1, N371, N378, ADD_22x22_fast_I126_Y_0, 
        N335, N332, N331, ADD_22x22_fast_I168_Y_0, \i_adj[10]_net_1 , 
        \i_adj[8]_net_1 , ADD_22x22_fast_I126_un1_Y_0, N379, 
        ADD_40x40_fast_I418_Y_0, ADD_22x22_fast_I177_Y_0, 
        \i_adj[19]_net_1 , \i_adj[17]_net_1 , ADD_22x22_fast_I179_Y_0, 
        \i_adj[21]_net_1 , ADD_22x22_fast_I130_Y_0, N386, 
        ADD_40x40_fast_I421_Y_0, N743, ADD_22x22_fast_I128_Y_0, N382, 
        N375, N374, ADD_22x22_fast_I127_Y_0, N380, N373, N372, 
        ADD_22x22_fast_I164_Y_0, \i_adj[4]_net_1 , \i_adj[6]_net_1 , 
        ADD_22x22_fast_I144_Y_2, ADD_22x22_fast_I144_un1_Y_0, N425, 
        ADD_22x22_fast_I144_Y_1, N369, N376, ADD_22x22_fast_I144_Y_0, 
        N333, N330, N329, ADD_22x22_fast_I143_Y_2, N367, 
        ADD_22x22_fast_I143_Y_1, N328, ADD_22x22_fast_I143_Y_0, N314, 
        ADD_22x22_fast_I142_Y_3, ADD_22x22_fast_I142_un1_Y_0, N421, 
        ADD_22x22_fast_I142_Y_2, N365, ADD_22x22_fast_I142_Y_1, N326, 
        ADD_22x22_fast_I142_Y_0, \i_adj[20]_net_1 , N317, 
        ADD_22x22_fast_I130_un1_Y_0, N387, \ireg[5]_net_1 , 
        \state[3]_net_1 , \ireg[23]_net_1 , \un1_next_sum_iv_0[4] , 
        \ireg[4]_net_1 , \ireg[20]_net_1 , \un1_next_sum_iv_0[22] , 
        \ireg[22]_net_1 , ADD_22x22_fast_I171_Y_0, \i_adj[11]_net_1 , 
        \i_adj[13]_net_1 , ADD_22x22_fast_I169_Y_0, \i_adj[9]_net_1 , 
        ADD_22x22_fast_I170_Y_0, \i_adj[12]_net_1 , 
        \un1_next_sum_iv_2[17] , \ireg[17]_net_1 , next_sum_0_sqmuxa, 
        \un1_next_sum_iv_0[17] , \un1_next_sum_iv_1[17] , \preg_m[17] , 
        \preg[17]_net_1 , next_sum_0_sqmuxa_2, next_sum_0_sqmuxa_1, 
        \un1_next_sum_iv_2[15] , \un3_next_sum_m[15] , 
        \un1_next_sum_iv_0[15] , \un1_next_sum_iv_1[15] , 
        \ireg[15]_net_1 , \preg_m[15] , \preg[15]_net_1 , 
        \un1_next_sum_iv_2[18] , \ireg[18]_net_1 , 
        \un1_next_sum_iv_0[18] , \un1_next_sum_iv_1[18] , \preg_m[18] , 
        \preg[18]_net_1 , \un1_next_sum_iv_2[12] , 
        \un24_next_sum_m[12] , \un3_next_sum_m[12] , 
        \un1_next_sum_iv_1[12] , \preg[12]_net_1 , \ireg_m[12] , 
        \ireg[16]_net_1 , \un1_next_sum_iv_0[16] , \preg_m[16] , 
        \preg[16]_net_1 , \ireg[11]_net_1 , \un1_next_sum_iv_0[11] , 
        \preg[11]_net_1 , \ireg_m[11] , \ireg[9]_net_1 , 
        \un1_next_sum_iv_0[9] , \preg[9]_net_1 , \ireg_m[9] , 
        \un1_next_sum_iv_2[13] , \un24_next_sum_m[13] , 
        \un3_next_sum_m[13] , \un1_next_sum_iv_1[13] , 
        \preg[13]_net_1 , \ireg_m[13] , \un1_next_sum_iv_2[8] , 
        \un24_next_sum_m[8] , \un3_next_sum_m[8] , 
        \un1_next_sum_iv_1[8] , \preg[8]_net_1 , \ireg_m[8] , 
        \un1_next_sum_iv_2[14] , \ireg[14]_net_1 , 
        \un1_next_sum_iv_0[14] , \un1_next_sum_iv_1[14] , \preg_m[14] , 
        \preg[14]_net_1 , \un1_next_sum_iv_2[7] , \un24_next_sum_m[7] , 
        \un3_next_sum_m[7] , \un1_next_sum_iv_1[7] , \preg[7]_net_1 , 
        \ireg_m[7] , \un1_next_sum_iv_2[6] , \un3_next_sum_m[6] , 
        \un1_next_sum_iv_0[6] , \un1_next_sum_iv_1[6] , 
        \preg[6]_net_1 , \ireg_m[6] , \un1_next_sum_iv_2[10] , 
        \un24_next_sum_m[10] , \un3_next_sum_m[10] , 
        \un1_next_sum_iv_1[10] , \preg[10]_net_1 , \ireg_m[10] , 
        ADD_22x22_fast_I128_un1_Y_0, N383, ADD_22x22_fast_I127_un1_Y_0, 
        N381, ADD_m8_i_1, ADD_m8_i_a4_0_0, \un1_next_sum_0_iv_1[25] , 
        \un3_next_sum_m[25] , ADD_22x22_fast_I129_Y_0, N384, N377, 
        ADD_22x22_fast_I165_Y_0, \i_adj[5]_net_1 , \i_adj[7]_net_1 , 
        ADD_22x22_fast_I129_un1_Y_0, N385, N266, N396, 
        ADD_22x22_fast_I162_Y_0, \i_adj[2]_net_1 , 
        ADD_22x22_fast_I163_Y_0, \i_adj[3]_net_1 , ADD_m8_i_a4_0_1, 
        ADD_m8_i_a4_0_0_0, ADD_m8_i_o4_1, 
        \un1_next_sum_0_sqmuxa_0_a4_1_0[0] , \state[4]_net_1 , 
        \state[5]_net_1 , ADD_m8_i_a4_2, N_232, \state[1]_net_1 , 
        N1031, I383_un1_Y, I340_un1_Y, N880, N745, N848, N1023, N819, 
        N597, N682, N1029, I382_un1_Y, I338_un1_Y, N878, N846, N1027, 
        I381_un1_Y, I336_un1_Y, N876, N823, N844, N1043, I286_un1_Y, 
        I348_un1_Y, N774, N790, N1091, N1040, N1088, N816, N734, N1049, 
        I290_un1_Y, I350_un1_Y, N778, N794, N1097, N1037, N1085, N1052, 
        I292_un1_Y, I351_un1_Y, N1100, N1035, I385_un1_Y, I344_un1_Y, 
        N884, N852, N1055, I294_un1_Y, N781, I352_un1_Y, N1103, N1046, 
        N1094, \next_ireg_3[25] , I120_un1_Y, \next_ireg_3[8] , N359, 
        \next_ireg_3[10] , N394, \next_ireg_3[11] , N531, 
        \next_ireg_3[16] , N422, I132_un1_Y, \next_ireg_3[7] , 
        \i_adj[1]_net_1 , \next_ireg_3[13] , N525, \next_ireg_3[20] , 
        \i_adj[14]_net_1 , N504, \next_ireg_3[21] , \i_adj[15]_net_1 , 
        N501, \next_ireg_3[22] , I126_un1_Y, \next_ireg_3[23] , 
        I124_un1_Y, \next_ireg_3[24] , N494, \next_ireg_3[19] , N507, 
        \next_ireg_3[18] , N510, \next_ireg_3[17] , N420, I131_un1_Y, 
        \next_ireg_3[15] , N424, I133_un1_Y, \next_ireg_3[14] , 
        I112_un1_Y, \next_ireg_3[12] , N528, \next_ireg_3[9] , 
        \ireg_m[25] , \un3_next_sum_m[24] , \ireg_m[24] , N680, N601, 
        N686, I353_un1_Y, N1106, N1058, I296_un1_Y, I378_un1_Y, N817, 
        N870, N838, N1021, I330_un1_Y, I380_un1_Y, N821, N874, N842, 
        N1025, I334_un1_Y, N882, N666, N850, N1033, N881, I143_un1_Y, 
        I122_un1_Y, N423, N407, N740, N478, N659, \next_sum[4] , 
        \next_sum[5] , \next_sum[6] , \next_sum[8] , \next_sum[9] , 
        \next_sum[10] , \next_sum[11] , \next_sum[12] , \next_sum[13] , 
        \next_sum[15] , \next_sum[16] , N1082, \next_sum[17] , N1079, 
        \next_sum[18] , N1076, \next_sum[19] , N1073, \next_sum[20] , 
        N1070, \next_sum[21] , N1067, \state[2]_net_1 , \next_sum[22] , 
        N1064, \next_sum[23] , N1061, \next_sum[24] , \next_sum[33] , 
        \next_sum[37] , N318, N388, N345, N342, N341, N293, N294, N346, 
        N389, N270, N272, N273, N278, N279, N282, N284, N285, N290, 
        N291, N296, N300, N343, N347, N351, N281, N352, N355, N356, 
        I87_un1_Y, N269, N344, N348, N354, N350, N390, N391, I86_un1_Y, 
        N340, N339, N299, N338, N337, N349, N336, N306, N287, N275, 
        \i_adj[0]_net_1 , N302, N305, N308, N311, N312, N334, N353, 
        N392, N357, N393, N358, I115_un1_Y, \next_ireg_3[6] , N795, 
        I308_un1_Y, I359_un1_Y, N705, N697, N729, N652, N649, N648, 
        N722, N645, N641, N721, N644, N640, N714, N637, N633, N713, 
        N636, N632, N709, N629, N628, N707, N630, N627, N626, N625, 
        N624, N703, I150_un1_Y, N622, N623, N617, N621, I144_un1_Y, 
        N616, N620, N495, N499, N498, N507_0, N511, N510_0, N519, 
        N525_0, N528_0, N532, N531_0, N535, N534, I66_un1_Y, N546, 
        N547, N538, N526, N520, N502, N496, N490, N487, N522, N486, 
        N541, N514, N517, N505, N653, N493, N704, N711, N634, N631, 
        N708, N710, N717, I358_un1_Y, N877, N875, N873, N869, 
        I320_un1_Y, N813, N814, N808, N807, N806, N805, N802, N801, 
        N797, I302_un1_Y, N789, I298_un1_Y, N799, N692, N739, N732, 
        I254_un1_Y, N731, N726, N733, N725, N724, I246_un1_Y, N723, 
        N728, N720, N718, N716, N700, N699, N696, N695, N688, N615, 
        N619, N693, I140_un1_Y, N613, N618, N540, N701, I70_un1_Y, 
        N639, N635, N647, N643, N651, N646, N642, N504_0, N501_0, N727, 
        N650, N654, N492, N489, N712, I230_un1_Y, N793, N719, N715, 
        N638, N516, N513, I242_un1_Y, \inf_abs1_5[0] , \inf_abs1_5[1] , 
        \inf_abs1_a_2[1] , \inf_abs1_5[2] , \inf_abs1_a_2[2] , 
        \inf_abs1_5[3] , \inf_abs1_a_2[3] , \inf_abs1_5[4] , 
        \inf_abs1_a_2[4] , \inf_abs1_5[5] , \inf_abs1_a_2[5] , 
        \inf_abs1_5[6] , \inf_abs1_a_2[6] , \inf_abs1_5[7] , 
        \inf_abs1_a_2[7] , \inf_abs1_5[8] , \inf_abs1_a_2[8] , 
        \inf_abs1_5[9] , \inf_abs1_a_2[9] , \inf_abs1_5[10] , 
        \inf_abs1_a_2[10] , \inf_abs1_5[11] , \inf_abs1_a_2[11] , 
        \inf_abs2_5[0] , \inf_abs2_5[1] , \inf_abs2_a_0[1] , 
        \inf_abs2_5[3] , \inf_abs2_a_0[3] , \inf_abs2_5[4] , 
        \inf_abs2_a_0[4] , \inf_abs2_5[5] , \inf_abs2_a_0[5] , 
        \inf_abs2_5[9] , \inf_abs2_a_0[9] , \inf_abs2_5[10] , 
        \inf_abs2_a_0[10] , \inf_abs2_5[11] , \inf_abs2_a_0[11] , 
        \inf_abs2_5[12] , \inf_abs2_a_0[12] , \inf_abs2_5[13] , 
        \inf_abs2_a_0[13] , \inf_abs2_5[17] , \inf_abs2_a_0[17] , 
        \inf_abs2_5[18] , \inf_abs2_a_0[18] , \inf_abs1_5[12] , 
        \inf_abs1_a_2[12] , \inf_abs2_5[19] , \inf_abs2_a_0[19] , 
        \inf_abs2_5[20] , \inf_abs2_a_0[20] , \inf_abs2_5[21] , 
        \inf_abs2_a_0[21] , \ireg[6]_net_1 , \ireg[7]_net_1 , 
        \ireg[8]_net_1 , \ireg[10]_net_1 , \ireg[12]_net_1 , 
        \ireg[13]_net_1 , \ireg[24]_net_1 , \ireg[25]_net_1 , 
        \inf_abs2_5[14] , \inf_abs2_a_0[14] , \inf_abs2_5[16] , 
        \inf_abs2_a_0[16] , \inf_abs2_5[8] , \inf_abs2_a_0[8] , N550, 
        N611, \next_sum[32] , \next_sum[28] , \next_sum[26] , 
        \next_sum[25] , N604, N605, N609, N606, N690, I212_un1_Y, 
        \next_sum[31] , N702, N694, I312_un1_Y, N815, I321_un1_Y, 
        I361_un1_Y, N483, N484, N656, \next_sum[27] , \next_sum[14] , 
        \next_sum[0] , N_228, \next_sum[2] , \next_sum[3] , N471, N481, 
        N741, I256_un1_Y, N662, N658, N480, N660, \state_ns[0] , N664, 
        I182_un1_Y, N735, N736, I250_un1_Y, N810, I306_un1_Y, 
        I318_un1_Y, N730, I184_un1_Y, N737, N738, N804, N812, 
        I259_un1_Y, N803, \next_sum[7] , \next_sum[1] , \next_sum[30] , 
        N607, N603, N610, N614, I252_un1_Y, I319_un1_Y, \next_sum[38] , 
        \next_sum[36] , \next_sum[35] , \next_sum[34] , \next_sum[29] , 
        \inf_abs2_5[15] , \inf_abs2_a_0[15] , \inf_abs2_5[7] , 
        \inf_abs2_a_0[7] , \inf_abs2_5[2] , \inf_abs2_a_0[2] , 
        \inf_abs2_5[6] , \inf_abs2_a_0[6] , \p_adj[0]_net_1 , 
        \p_adj[1]_net_1 , \p_adj[2]_net_1 , \p_adj[3]_net_1 , 
        \p_adj[4]_net_1 , \p_adj[5]_net_1 , \p_adj[6]_net_1 , 
        \p_adj[7]_net_1 , \p_adj[8]_net_1 , \p_adj[9]_net_1 , 
        \p_adj[10]_net_1 , \p_adj[11]_net_1 , \p_adj[12]_net_1 , N_6, 
        \DWACT_FINC_E[28] , \DWACT_FINC_E[13] , \DWACT_FINC_E[15] , 
        N_7, \DWACT_FINC_E[14] , N_8, \DWACT_FINC_E[9] , 
        \DWACT_FINC_E[12] , N_9, \DWACT_FINC_E[10] , \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[5] , N_10_0, \DWACT_FINC_E[11] , N_11, N_12_0, 
        N_13, \DWACT_FINC_E[8] , N_14, N_16, N_17, \DWACT_FINC_E[3] , 
        N_19, N_20, N_21, \DWACT_FINC_E[1] , N_22, N_24, N_3, 
        \DWACT_FINC_E_0[2] , \DWACT_FINC_E_0[5] , N_4, 
        \DWACT_FINC_E_0[3] , N_6_0, N_7_0, N_8_0, \DWACT_FINC_E_0[1] , 
        N_9_0, N_11_0, GND, VCC;
    
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I312_un1_Y (.A(N815), .B(N800), 
        .Y(I312_un1_Y));
    DFN1E1C0 \sumreg[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(sum_39));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I77_Y (.A(sum_19), .B(
        \un1_next_sum[19] ), .C(N532), .Y(N627));
    XA1B \state_RNIJBKS5A[2]  (.A(N1021), .B(ADD_40x40_fast_I457_Y_0), 
        .C(\state[2]_net_1 ), .Y(\next_sum[39] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I19_G0N (.A(\un1_next_sum[19] )
        , .B(sum_19), .Y(N528_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I14_P0N (.A(\un1_next_sum[14] ), 
        .B(sum_14), .Y(N514));
    NOR3B \preg_RNIPEAK[12]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[12]_net_1 ), .Y(\un24_next_sum_m[12] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I46_Y (.A(\sumreg[35]_net_1 ), 
        .B(\sumreg[34]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N596)
        );
    XA1B \sumreg_RNO[10]  (.A(N1100), .B(ADD_40x40_fast_I428_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[10] ));
    MX2 \p_adj_RNO[2]  (.A(sr_new[2]), .B(\inf_abs1_a_2[2] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[2] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I336_un1_Y (.A(N844), .B(N875), 
        .Y(I336_un1_Y));
    XA1B \sumreg_RNO[11]  (.A(N1097), .B(ADD_40x40_fast_I429_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[11] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_0 (.A(N333), .B(N330), .C(
        N329), .Y(ADD_22x22_fast_I144_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I241_Y (.A(N718), .B(N726), .Y(
        N800));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I114_Y (.A(N471), .B(
        \un1_next_sum[0] ), .C(sum_1_d0), .Y(N664));
    DFN1E1C0 \i_adj[19]  (.D(\inf_abs2_5[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[19]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I113_Y (.A(N389), .B(N396), .C(
        N388), .Y(N525));
    DFN1E1C0 \sumreg[23]  (.D(\next_sum[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(sum_23));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I290_un1_Y (.A(N793), .B(N778), 
        .Y(I290_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I128_un1_Y_0 (.A(N383), .B(N375)
        , .Y(ADD_22x22_fast_I128_un1_Y_0));
    NOR3B inf_abs1_a_2_I_19 (.A(\DWACT_FINC_E_0[2] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[6]), .Y(N_7_0));
    OA1 next_ireg_3_0_ADD_22x22_fast_I33_Y (.A(\i_adj[12]_net_1 ), .B(
        \i_adj[14]_net_1 ), .C(N300), .Y(N338));
    NOR3B \ireg_RNIBUL41[8]  (.A(\state[3]_net_1 ), .B(\ireg[8]_net_1 )
        , .C(integral_1_0), .Y(\ireg_m[8] ));
    AND3 inf_abs2_a_0_I_30 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E_0[6] ));
    MX2 \i_adj_RNO[5]  (.A(integral[11]), .B(\inf_abs2_a_0[5] ), .S(
        integral_0_0), .Y(\inf_abs2_5[5] ));
    AO1 \ireg_RNI5S191[15]  (.A(\ireg[15]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[15] ), .Y(
        \un1_next_sum_iv_1[15] ));
    XA1 \ireg_RNI57LQ[22]  (.A(integral_0_0), .B(\ireg[22]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[22] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I304_Y (.A(N807), .B(N792), .C(
        N791), .Y(N875));
    DFN1E1C0 \sumreg[38]  (.D(\next_sum[38] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[38]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I126_un1_Y_0 (.A(N371), .B(N379)
        , .Y(ADD_22x22_fast_I126_un1_Y_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I361_Y (.A(N799), .B(I312_un1_Y), 
        .C(I361_un1_Y), .Y(N1082));
    DFN1E1C0 \sumreg[5]  (.D(\next_sum[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_5));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I248_Y (.A(N733), .B(N726), .C(
        N725), .Y(N807));
    DFN1E1C0 \sumreg[20]  (.D(\next_sum[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(sum_20));
    AO1 next_ireg_3_0_ADD_22x22_fast_I128_Y (.A(
        ADD_22x22_fast_I128_un1_Y_0), .B(N528), .C(
        ADD_22x22_fast_I128_Y_0), .Y(N504));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I150_un1_Y (.A(N626), .B(N623), 
        .Y(I150_un1_Y));
    NOR2 inf_abs2_a_0_I_57 (.A(integral[24]), .B(integral[25]), .Y(
        \DWACT_FINC_E[14] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I378_Y_1 (.A(
        ADD_40x40_fast_I378_Y_0), .B(N594), .Y(ADD_40x40_fast_I378_Y_1)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I347_Y_0 (.A(N787), .B(N772), .C(
        N771), .Y(ADD_40x40_fast_I347_Y_0));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I52_Y (.A(\sumreg[31]_net_1 ), 
        .B(\sumreg[32]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N602)
        );
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I199_Y (.A(
        ADD_40x40_fast_I199_Y_0), .B(N684), .Y(N758));
    AO1 \ireg_RNI90291[17]  (.A(\ireg[17]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[17] ), .Y(
        \un1_next_sum_iv_1[17] ));
    DFN1E1C0 \sumreg[13]  (.D(\next_sum[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_13));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I354_Y (.A(N870), .B(N817), .C(
        N869), .Y(N1061));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I214_Y (.A(N699), .B(N692), .C(
        N691), .Y(N773));
    OA1 next_ireg_3_0_ADD_22x22_fast_I21_Y (.A(\i_adj[18]_net_1 ), .B(
        \i_adj[20]_net_1 ), .C(N318), .Y(N326));
    NOR3B \ireg_RNIPK7P[24]  (.A(\state[3]_net_1 ), .B(
        \ireg[24]_net_1 ), .C(integral_1_0), .Y(\ireg_m[24] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I353_un1_Y_0 (.A(N800), .B(
        N784), .Y(ADD_40x40_fast_I353_un1_Y_0));
    DFN1E1C0 \i_adj[2]  (.D(\inf_abs2_5[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[2]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I225_Y (.A(N702), .B(N710), .Y(
        N784));
    NOR3A inf_abs1_a_2_I_13 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .C(
        sr_new[4]), .Y(N_9_0));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I436_Y_0 (.A(sum_18), .B(
        \un1_next_sum[18] ), .Y(ADD_40x40_fast_I436_Y_0));
    DFN1E1C0 \sumreg[27]  (.D(\next_sum[27] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[27]_net_1 ));
    DFN1E1C0 \sumreg[10]  (.D(\next_sum[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_10));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I381_Y_2 (.A(N760), .B(N775), .C(
        ADD_40x40_fast_I381_Y_1), .Y(ADD_40x40_fast_I381_Y_2));
    NOR2 \state_RNI19LH[4]  (.A(\state[4]_net_1 ), .B(\state[5]_net_1 )
        , .Y(\un1_next_sum_0_sqmuxa_0_a4_1_0[0] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I15_P0N (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(N312));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I444_Y_0 (.A(
        \sumreg[26]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I444_Y_0));
    XA1B \sumreg_RNO[22]  (.A(N1064), .B(ADD_40x40_fast_I440_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[22] ));
    OR3 \ireg_RNIUMS52[12]  (.A(\un24_next_sum_m[12] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[12] ), .Y(
        \un1_next_sum_iv_2[12] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I171_Y (.A(N647), .B(N643), .Y(
        N724));
    OR2 \un1_next_sum_iv[21]  (.A(N_228_1), .B(
        \un1_next_sum_iv_0[21]_net_1 ), .Y(\un1_next_sum[21] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I11_P0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(N300));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I443_Y_0 (.A(
        \sumreg[25]_net_1 ), .B(\un1_next_sum_0_iv[25] ), .Y(
        ADD_40x40_fast_I443_Y_0));
    AND2 inf_abs2_a_0_I_44 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E[9] ), .Y(\DWACT_FINC_E[10] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I18_P0N (.A(\un1_next_sum[18] ), 
        .B(sum_18), .Y(N526));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I306_un1_Y (.A(N727), .B(
        I250_un1_Y), .C(N794), .Y(I306_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I166_Y (.A(N642), .B(N639), .C(
        N638), .Y(N719));
    OR2 \preg_RNI31Q64[8]  (.A(\un1_next_sum_iv_2[8] ), .B(
        \un1_next_sum_iv_1[8] ), .Y(\un1_next_sum[8] ));
    AX1D next_ireg_3_0_ADD_22x22_fast_I168_Y (.A(N386), .B(I112_un1_Y), 
        .C(ADD_22x22_fast_I168_Y_0), .Y(\next_ireg_3[14] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I10_G0N (.A(\un1_next_sum[10] )
        , .B(sum_10), .Y(N501_0));
    XNOR2 inf_abs1_a_2_I_28 (.A(sr_new[10]), .B(N_4), .Y(
        \inf_abs1_a_2[10] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I18_G0N (.A(\un1_next_sum[18] )
        , .B(sum_18), .Y(N525_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I338_un1_Y (.A(N846), .B(N877), 
        .Y(I338_un1_Y));
    DFN1E1C0 \p_adj[4]  (.D(\inf_abs1_5[4] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[4]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_2 (.A(
        ADD_22x22_fast_I144_un1_Y_0), .B(N425), .C(
        ADD_22x22_fast_I144_Y_1), .Y(ADD_22x22_fast_I144_Y_2));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I358_Y (.A(I358_un1_Y), .B(N877), 
        .Y(N1073));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I7_G0N (.A(\i_adj[7]_net_1 ), 
        .B(\i_adj[9]_net_1 ), .Y(N287));
    XNOR2 inf_abs2_a_0_I_20 (.A(integral[13]), .B(N_20), .Y(
        \inf_abs2_a_0[7] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I424_Y_0 (.A(sum_6), .B(
        \un1_next_sum[6] ), .Y(ADD_40x40_fast_I424_Y_0));
    DFN1E1C0 \sumreg[17]  (.D(\next_sum[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_17));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I257_Y_1 (.A(N475), .B(N472), 
        .C(N661), .Y(ADD_40x40_fast_I257_Y_1));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I321_Y (.A(I321_un1_Y), .B(N815), 
        .Y(N1106));
    DFN1C0 \state[6]  (.D(\state_2[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[6]_net_1 ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I423_Y_0 (.A(N_228_1), .B(
        \un1_next_sum_iv_0[5] ), .C(sum_5), .Y(ADD_40x40_fast_I423_Y_0)
        );
    AND3 inf_abs1_a_2_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[5] ), .Y(
        \DWACT_FINC_E[6] ));
    DFN1E1C0 \sumreg[35]  (.D(\next_sum[35] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[35]_net_1 ));
    MX2 \i_adj_RNO[13]  (.A(integral[19]), .B(\inf_abs2_a_0[13] ), .S(
        integral_1_0), .Y(\inf_abs2_5[13] ));
    DFN1E1C0 \sumreg[4]  (.D(\next_sum[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_4));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I87_un1_Y (.A(N358), .B(N266), 
        .Y(I87_un1_Y));
    XA1B \sumreg_RNO[38]  (.A(N1023), .B(ADD_40x40_fast_I456_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[38] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I160_Y (.A(N636), .B(N633), .C(
        N632), .Y(N713));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I232_Y (.A(N717), .B(N710), .C(
        N709), .Y(N791));
    NOR2 inf_abs2_a_0_I_6 (.A(integral[6]), .B(integral[7]), .Y(N_25));
    NOR3B inf_abs2_a_0_I_45 (.A(\DWACT_FINC_E[10] ), .B(
        \DWACT_FINC_E_0[6] ), .C(integral[21]), .Y(N_11));
    NOR3 inf_abs1_a_2_I_29 (.A(sr_new[7]), .B(sr_new[6]), .C(sr_new[8])
        , .Y(\DWACT_FINC_E_0[5] ));
    NOR2A \state_RNIHR1J_0[3]  (.A(\state[3]_net_1 ), .B(integral[25]), 
        .Y(next_sum_1_sqmuxa));
    NOR2B \ireg_RNIACOK[25]  (.A(\ireg[25]_net_1 ), .B(
        next_sum_0_sqmuxa), .Y(\ireg_m[25] ));
    MX2 \p_adj_RNO[1]  (.A(sr_new[1]), .B(\inf_abs1_a_2[1] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[1] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I382_un1_Y (.A(N878), .B(N743), 
        .C(N846), .Y(I382_un1_Y));
    OR2 \un1_next_sum_iv_0[21]  (.A(\un3_next_sum_m[21] ), .B(
        \ireg_m[21] ), .Y(\un1_next_sum_iv_0[21]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I252_un1_Y (.A(N737), .B(N730), 
        .Y(I252_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I53_Y (.A(N270), .B(N273), .Y(
        N358));
    AO1 next_ireg_3_0_ADD_22x22_fast_I30_Y (.A(N302), .B(N306), .C(
        N305), .Y(N335));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I124_un1_Y (.A(N377), .B(N369), 
        .C(N424), .Y(I124_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I330_un1_Y (.A(N838), .B(N869), 
        .Y(I330_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I237_Y (.A(N722), .B(N714), .Y(
        N796));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I12_G0N (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[12]_net_1 ), .Y(N302));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I11_G0N (.A(\i_adj[13]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(N299));
    OR2 \ireg_RNIN7293[18]  (.A(\un1_next_sum_iv_2[18] ), .B(
        \un1_next_sum_iv_1[18] ), .Y(\un1_next_sum[18] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I58_Y (.A(\sumreg[28]_net_1 ), 
        .B(\sumreg[29]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N608)
        );
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I257_Y (.A(
        ADD_40x40_fast_I257_Y_1), .B(N734), .Y(N816));
    NOR2B \state_RNIHR1J[3]  (.A(\state[3]_net_1 ), .B(integral[25]), 
        .Y(next_sum_0_sqmuxa));
    OA1 next_ireg_3_0_ADD_22x22_fast_I35_Y (.A(\i_adj[12]_net_1 ), .B(
        \i_adj[10]_net_1 ), .C(N300), .Y(N340));
    NOR2B un1_sumreg_0_0_ADD_m8_i_a4_0_0 (.A(sum_0_d0), .B(sum_1_d0), 
        .Y(ADD_m8_i_a4_0_0_0));
    DFN1E1C0 \sumreg[7]  (.D(\next_sum[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_7));
    DFN1E1C0 \ireg[12]  (.D(\next_ireg_3[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[12]_net_1 ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I176_Y_0 (.A(\i_adj[18]_net_1 ), 
        .B(\i_adj[16]_net_1 ), .Y(ADD_22x22_fast_I176_Y_0));
    NOR2A inf_abs2_a_0_I_11 (.A(\DWACT_FINC_E_0[0] ), .B(integral[9]), 
        .Y(N_23));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I166_Y (.A(\i_adj[6]_net_1 ), .B(
        \i_adj[8]_net_1 ), .C(N528), .Y(\next_ireg_3[12] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I67_Y (.A(\sumreg[24]_net_1 ), 
        .B(\un1_next_sum[24] ), .C(N547), .Y(N617));
    AO1 next_ireg_3_0_ADD_22x22_fast_I38_Y (.A(N290), .B(N294), .C(
        N293), .Y(N343));
    XNOR2 inf_abs2_a_0_I_46 (.A(integral[22]), .B(N_11), .Y(
        \inf_abs2_a_0[16] ));
    XOR2 inf_abs1_a_2_I_5 (.A(sr_new[0]), .B(sr_new[1]), .Y(
        \inf_abs1_a_2[1] ));
    XNOR2 inf_abs1_a_2_I_23 (.A(sr_new[8]), .B(N_6_0), .Y(
        \inf_abs1_a_2[8] ));
    OR3 \state_RNIFG0J1_0[4]  (.A(next_sum_1_sqmuxa_2), .B(
        next_sum_1_sqmuxa_1), .C(next_sum_1_sqmuxa), .Y(
        \un1_next_sum_1_iv[26] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I310_Y (.A(N813), .B(N798), .C(
        N797), .Y(N881));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I308_un1_Y (.A(N729), .B(
        I252_un1_Y), .C(N796), .Y(I308_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I169_Y (.A(N645), .B(N641), .Y(
        N722));
    AO1A \preg_RNI0O8B1[18]  (.A(\preg[18]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[18] ));
    DFN1C0 \state[2]  (.D(\state[1]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[2]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I245_Y (.A(N730), .B(N722), .Y(
        N804));
    DFN1E1C0 \i_adj[15]  (.D(\inf_abs2_5[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[15]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I349_Y_0 (.A(N791), .B(N776), .C(
        N775), .Y(ADD_40x40_fast_I349_Y_0));
    OA1 next_ireg_3_0_ADD_22x22_fast_I41_Y (.A(\i_adj[9]_net_1 ), .B(
        \i_adj[7]_net_1 ), .C(N291), .Y(N346));
    DFN1E1C0 \i_adj[20]  (.D(\inf_abs2_5[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[20]_net_1 ));
    XNOR2 inf_abs2_a_0_I_37 (.A(integral[19]), .B(N_14), .Y(
        \inf_abs2_a_0[13] ));
    MX2 \i_adj_RNO[12]  (.A(integral[18]), .B(\inf_abs2_a_0[12] ), .S(
        integral_1_0), .Y(\inf_abs2_5[12] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I53_Y (.A(\sumreg[32]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N603)
        );
    OR2 next_ireg_3_0_ADD_22x22_fast_I86_Y (.A(I86_un1_Y), .B(N355), 
        .Y(N394));
    AX1D next_ireg_3_0_ADD_22x22_fast_I170_Y (.A(N422), .B(I132_un1_Y), 
        .C(ADD_22x22_fast_I170_Y_0), .Y(\next_ireg_3[16] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I144_Y_1 (.A(N369), .B(N376), .C(
        ADD_22x22_fast_I144_Y_0), .Y(ADD_22x22_fast_I144_Y_1));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I4_P0N (.A(\un1_next_sum[4] ), 
        .B(sum_4), .Y(N484));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I213_Y (.A(N690), .B(N698), .Y(
        N772));
    DFN1E1C0 \p_adj[10]  (.D(\inf_abs1_5[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[10]_net_1 ));
    DFN1E1C0 \p_adj[5]  (.D(\inf_abs1_5[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[5]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I164_Y (.A(N640), .B(N637), .C(
        N636), .Y(N717));
    DFN1E1C0 \sumreg[36]  (.D(\next_sum[36] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[36]_net_1 ));
    NOR3B \ireg_RNI56KQ[13]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[13]_net_1 ), .Y(\un3_next_sum_m[13] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I56_Y (.A(\sumreg[30]_net_1 ), 
        .B(\sumreg[29]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N606)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I172_Y (.A(N648), .B(N645), .C(
        N644), .Y(N725));
    NOR2B \p_adj_RNO[12]  (.A(\inf_abs1_a_2[12] ), .B(sr_new[12]), .Y(
        \inf_abs1_5[12] ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I126_un1_Y (.A(N386), .B(
        I112_un1_Y), .C(ADD_22x22_fast_I126_un1_Y_0), .Y(I126_un1_Y));
    DFN1E1C0 \p_adj[0]  (.D(\inf_abs1_5[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[0]_net_1 ));
    AND3 inf_abs2_a_0_I_51 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[28] ));
    DFN1E1C0 \sumreg[9]  (.D(\next_sum[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_9));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I181_Y (.A(N487), .B(N484), .C(
        N653), .Y(N734));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I216_Y (.A(N701), .B(N694), .C(
        N693), .Y(N775));
    OA1 un1_sumreg_0_0_ADD_m8_i_a4 (.A(N_232), .B(ADD_m8_i_o4_1), .C(
        next_sum_0_sqmuxa), .Y(ADD_m8_i_a4_2));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I4_G0N (.A(\un1_next_sum[4] ), 
        .B(sum_4), .Y(N483));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I317_Y (.A(N808), .B(N823), .C(
        N807), .Y(N1094));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I129_Y (.A(N601), .B(N605), .Y(
        N682));
    OR3 \preg_RNIADKC2[8]  (.A(\un24_next_sum_m[8] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[8] ), .Y(
        \un1_next_sum_iv_2[8] ));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I50_Y (.A(N272), .B(
        \i_adj[3]_net_1 ), .C(\i_adj[5]_net_1 ), .Y(N355));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I144_un1_Y_0 (.A(N377), .B(N369)
        , .C(N266), .Y(ADD_22x22_fast_I144_un1_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I34_Y (.A(N296), .B(N300), .C(
        N299), .Y(N339));
    OR3 \ireg_RNIQIS52[10]  (.A(\un24_next_sum_m[10] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[10] ), .Y(
        \un1_next_sum_iv_2[10] ));
    DFN1E1C0 \sumreg[31]  (.D(\next_sum[31] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[31]_net_1 ));
    DFN1E1C0 \sumreg[2]  (.D(\next_sum[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_2_d0));
    DFN1E1C0 \i_adj[7]  (.D(\inf_abs2_5[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[7]_net_1 ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I383_Y (.A(
        ADD_40x40_fast_I383_Y_1), .B(I383_un1_Y), .C(I340_un1_Y), .Y(
        N1031));
    MX2 \i_adj_RNO[8]  (.A(integral[14]), .B(\inf_abs2_a_0[8] ), .S(
        integral_0_0), .Y(\inf_abs2_5[8] ));
    NOR3B \ireg_RNIQJ601[7]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[7]_net_1 ), .Y(\un3_next_sum_m[7] ));
    AO1A \ireg_RNIUMVV1[11]  (.A(\ireg[11]_net_1 ), .B(
        next_sum_0_sqmuxa), .C(\un1_next_sum_iv_0[11] ), .Y(
        \un1_next_sum_iv_2[11] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I9_P0N (.A(
        \un1_next_sum_iv_1[9] ), .B(\un1_next_sum_iv_2[9] ), .C(sum_9), 
        .Y(N499));
    NOR3A inf_abs2_a_0_I_27 (.A(\DWACT_FINC_E_0[4] ), .B(integral[14]), 
        .C(integral[15]), .Y(N_17));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I10_G0N (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[12]_net_1 ), .Y(N296));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I351_un1_Y_0 (.A(N706), .B(
        N698), .C(N796), .Y(ADD_40x40_fast_I351_un1_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I108_Y (.A(N390), .B(N383), .C(
        N382), .Y(N422));
    MX2 \p_adj_RNO[3]  (.A(sr_new[3]), .B(\inf_abs1_a_2[3] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[3] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I435_Y_0 (.A(sum_17), .B(
        \un1_next_sum[17] ), .Y(ADD_40x40_fast_I435_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I146_Y (.A(N622), .B(N619), .C(
        N618), .Y(N699));
    AND3 inf_abs2_a_0_I_48 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[11] ), .Y(N_10_0));
    OA1A un1_sumreg_0_0_ADD_40x40_fast_I197_Y_0 (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[36]_net_1 ), .C(N583), .Y(
        ADD_40x40_fast_I197_Y_0));
    DFN1E1C0 \preg[16]  (.D(\p_adj[10]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[16]_net_1 ));
    NOR3B \ireg_RNICVL41[9]  (.A(\state[3]_net_1 ), .B(\ireg[9]_net_1 )
        , .C(integral_1_0), .Y(\ireg_m[9] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I135_Y (.A(N607), .B(N611), .Y(
        N688));
    DFN1E1C0 \preg[17]  (.D(\p_adj[11]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[17]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I9_G0N (.A(\i_adj[9]_net_1 ), 
        .B(\i_adj[11]_net_1 ), .Y(N293));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I155_Y (.A(N627), .B(N631), .Y(
        N708));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I122_un1_Y (.A(N407), .B(N422), 
        .Y(I122_un1_Y));
    OR2 next_ireg_3_0_ADD_22x22_fast_I5_P0N (.A(\i_adj[7]_net_1 ), .B(
        \i_adj[5]_net_1 ), .Y(N282));
    DFN1E1C0 \i_adj[8]  (.D(\inf_abs2_5[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[8]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I94_Y (.A(N501_0), .B(N505), .C(
        N504_0), .Y(N644));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I73_Y (.A(N346), .B(N342), .Y(
        N381));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I174_Y (.A(\i_adj[16]_net_1 ), 
        .B(\i_adj[14]_net_1 ), .C(N504), .Y(\next_ireg_3[20] ));
    DFN1E1C0 \i_adj[17]  (.D(\inf_abs2_5[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[17]_net_1 ));
    AO1A \preg_RNIPG8B1[11]  (.A(\preg[11]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[11] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I140_Y (.A(I140_un1_Y), .B(N612), 
        .Y(N693));
    MX2 \i_adj_RNO[3]  (.A(integral[9]), .B(\inf_abs2_a_0[3] ), .S(
        integral_0_0), .Y(\inf_abs2_5[3] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I74_Y (.A(N531_0), .B(N535), .C(
        N534), .Y(N624));
    XNOR2 inf_abs2_a_0_I_49 (.A(integral[23]), .B(N_10_0), .Y(
        \inf_abs2_a_0[17] ));
    OR2 \ireg_RNI4TS52[15]  (.A(\un3_next_sum_m[15] ), .B(
        \un1_next_sum_iv_0[15] ), .Y(\un1_next_sum_iv_2[15] ));
    XNOR2 inf_abs2_a_0_I_12 (.A(integral[10]), .B(N_23), .Y(
        \inf_abs2_a_0[4] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I319_Y (.A(N729), .B(I252_un1_Y), 
        .C(I319_un1_Y), .Y(N1100));
    XA1B \sumreg_RNO[18]  (.A(N1076), .B(ADD_40x40_fast_I436_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[18] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I306_Y (.A(I306_un1_Y), .B(N793), 
        .Y(N877));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I224_Y (.A(N709), .B(N702), .C(
        N701), .Y(N783));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I209_Y (.A(N686), .B(N694), .Y(
        N768));
    OR2 \state_RNIUKUV[5]  (.A(next_sum_0_sqmuxa_1), .B(
        next_sum_0_sqmuxa_2), .Y(N_228_1));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I383_Y_0 (.A(N608), .B(N612), .C(
        N681), .Y(ADD_40x40_fast_I383_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I17_G0N (.A(\un1_next_sum[17] )
        , .B(sum_17), .Y(N522));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I356_Y (.A(N874), .B(N821), .C(
        N873), .Y(N1067));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I239_Y (.A(N716), .B(N724), .Y(
        N798));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I259_Y (.A(I259_un1_Y), .B(N737), 
        .Y(N819));
    NOR3B \ireg_RNI59QU[12]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[12]_net_1 ), .C(integral_1_0), .Y(\ireg_m[12] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I106_Y (.A(N388), .B(N381), .C(
        N380), .Y(N420));
    NOR2B \i_adj_RNO[21]  (.A(\inf_abs2_a_0[21] ), .B(integral[25]), 
        .Y(\inf_abs2_5[21] ));
    DFN1E1C0 \sumreg[6]  (.D(\next_sum[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_6));
    DFN1E1C0 \sumreg[0]  (.D(\next_sum[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_0_d0));
    DFN1E1C0 \preg[15]  (.D(\p_adj[9]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[15]_net_1 ));
    DFN1E1C0 \i_adj[10]  (.D(\inf_abs2_5[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[10]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I144_un1_Y (.A(N620), .B(N617), 
        .Y(I144_un1_Y));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I452_Y_0 (.A(
        \sumreg[34]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I452_Y_0));
    DFN1E1C0 \ireg[24]  (.D(\next_ireg_3[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[24]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I271_Y (.A(N758), .B(N774), .Y(
        N842));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I351_un1_Y (.A(
        ADD_40x40_fast_I351_un1_Y_0), .B(N1100), .Y(I351_un1_Y));
    XNOR2 inf_abs2_a_0_I_43 (.A(integral[21]), .B(N_12_0), .Y(
        \inf_abs2_a_0[15] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I69_Y (.A(N338), .B(N342), .Y(
        N377));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I385_Y (.A(I385_un1_Y), .B(
        ADD_40x40_fast_I385_Y_1), .C(I344_un1_Y), .Y(N1035));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I184_un1_Y (.A(N487), .B(N484), 
        .C(N660), .Y(I184_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I149_Y (.A(N625), .B(N621), .Y(
        N702));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I67_Y (.A(N336), .B(N340), .Y(
        N375));
    OR2 next_ireg_3_0_ADD_22x22_fast_I54_Y (.A(I87_un1_Y), .B(N269), 
        .Y(N359));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I378_Y_2 (.A(N598), .B(N602), .C(
        ADD_40x40_fast_I378_Y_1), .Y(ADD_40x40_fast_I378_Y_2));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I360_Y (.A(N882), .B(N666), .C(
        N881), .Y(N1079));
    MX2 \p_adj_RNO[0]  (.A(sr_new[0]), .B(sr_new[0]), .S(sr_new_0_0), 
        .Y(\inf_abs1_5[0] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I384_Y_0 (.A(N691), .B(N684), .C(
        N683), .Y(ADD_40x40_fast_I384_Y_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I182_Y (.A(I182_un1_Y), .B(N654), 
        .Y(N735));
    OR2 \un1_next_sum_iv_0[19]  (.A(\un3_next_sum_m[19] ), .B(
        \ireg_m[19] ), .Y(\un1_next_sum_iv_0[19]_net_1 ));
    AND3 inf_abs2_a_0_I_52 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[12] ), .Y(N_9));
    NOR3A inf_abs2_a_0_I_31 (.A(\DWACT_FINC_E_0[6] ), .B(integral[15]), 
        .C(integral[16]), .Y(N_16));
    OR2 \preg_RNIK61P3[10]  (.A(\un1_next_sum_iv_2[10] ), .B(
        \un1_next_sum_iv_1[10] ), .Y(\un1_next_sum[10] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I163_Y (.A(N639), .B(N635), .Y(
        N716));
    AO1 next_ireg_3_0_ADD_22x22_fast_I110_Y (.A(N392), .B(N385), .C(
        N384), .Y(N424));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I197_Y (.A(N597), .B(
        ADD_40x40_fast_I197_Y_0), .C(N682), .Y(N756));
    NOR2B \state_RNITH09[5]  (.A(\state[5]_net_1 ), .B(sr_new[12]), .Y(
        next_sum_0_sqmuxa_2));
    DFN1E1C0 \i_adj[18]  (.D(\inf_abs2_5[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[18]_net_1 ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I91_Y (.A(sum_12), .B(
        \un1_next_sum[12] ), .C(N511), .Y(N641));
    NOR3B \preg_RNINCAK[10]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[10]_net_1 ), .Y(\un24_next_sum_m[10] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I93_Y (.A(N367), .B(N375), .Y(
        N407));
    OR2A un1_sumreg_0_0_ADD_40x40_fast_I25_P0N (.A(
        \un1_next_sum_0_iv[25] ), .B(\sumreg[25]_net_1 ), .Y(N547));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I144_Y (.A(I144_un1_Y), .B(N616), 
        .Y(N697));
    OR2 \state_RNIH6RR1[4]  (.A(N_228_1), .B(N_232), .Y(N_228));
    MX2 \i_adj_RNO[16]  (.A(integral[22]), .B(\inf_abs2_a_0[16] ), .S(
        integral_1_0), .Y(\inf_abs2_5[16] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I71_Y (.A(N541), .B(N538), .Y(
        N621));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I95_Y (.A(N505), .B(N502), .Y(
        N645));
    OR2 next_ireg_3_0_ADD_22x22_fast_I13_P0N (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[13]_net_1 ), .Y(N306));
    AND2 un1_sumreg_0_0_ADD_40x40_fast_I195_Y_1 (.A(N595), .B(
        ADD_40x40_fast_I195_Y_0), .Y(ADD_40x40_fast_I195_Y_1));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I319_un1_Y (.A(N812), .B(N745), 
        .Y(I319_un1_Y));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I161_Y (.A(\i_adj[3]_net_1 ), .B(
        \i_adj[1]_net_1 ), .C(N266), .Y(\next_ireg_3[7] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I70_Y (.A(N343), .B(N340), .C(
        N339), .Y(N378));
    AO1A \ireg_RNICFKC2[9]  (.A(\ireg[9]_net_1 ), .B(next_sum_0_sqmuxa)
        , .C(\un1_next_sum_iv_0[9] ), .Y(\un1_next_sum_iv_2[9] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I75_Y (.A(N532), .B(N535), .Y(
        N625));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I168_Y (.A(N644), .B(N641), .C(
        N640), .Y(N721));
    MX2 \p_adj_RNO[6]  (.A(sr_new[6]), .B(\inf_abs1_a_2[6] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[6] ));
    OR3 \ireg_RNIVM1O2[24]  (.A(\un3_next_sum_m[24] ), .B(\ireg_m[24] )
        , .C(N_228_1), .Y(\un1_next_sum[24] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I379_Y_3 (.A(N756), .B(N771), .C(
        ADD_40x40_fast_I379_Y_2), .Y(ADD_40x40_fast_I379_Y_3));
    NOR2B \state_RNIJHSR[4]  (.A(\un1_next_sum_0_sqmuxa_0_a4_1_0[0] ), 
        .B(integral[25]), .Y(N_232));
    AO1A \preg_RNIVM8B1[17]  (.A(\preg[17]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[17] ));
    NOR2B \preg_RNIRGAK[14]  (.A(\preg[14]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[14] ));
    MX2 \i_adj_RNO[1]  (.A(integral[7]), .B(\inf_abs2_a_0[1] ), .S(
        integral_0_0), .Y(\inf_abs2_5[1] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I75_Y (.A(N344), .B(N348), .Y(
        N383));
    GND GND_i (.Y(GND));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I143_Y_0 (.A(\i_adj[17]_net_1 ), 
        .B(\i_adj[19]_net_1 ), .C(N314), .Y(ADD_22x22_fast_I143_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I244_Y (.A(N729), .B(N722), .C(
        N721), .Y(N803));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I314_Y (.A(N802), .B(N817), .C(
        N801), .Y(N1085));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I320_Y (.A(I320_un1_Y), .B(N813), 
        .Y(N1103));
    AO1A \preg_RNITK8B1[15]  (.A(\preg[15]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[15] ));
    MX2 \p_adj_RNO[5]  (.A(sr_new[5]), .B(\inf_abs1_a_2[5] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[5] ));
    OR2 \preg_RNI0J1P3[13]  (.A(\un1_next_sum_iv_2[13] ), .B(
        \un1_next_sum_iv_1[13] ), .Y(\un1_next_sum[13] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I378_Y_3 (.A(N754), .B(N769), .C(
        ADD_40x40_fast_I378_Y_2), .Y(ADD_40x40_fast_I378_Y_3));
    DFN1C0 \state[5]  (.D(\state[4]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[5]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I78_Y (.A(N351), .B(N348), .C(
        N347), .Y(N386));
    AO1A \ireg_RNIC5002[18]  (.A(\ireg[18]_net_1 ), .B(
        next_sum_0_sqmuxa), .C(\un1_next_sum_iv_0[18] ), .Y(
        \un1_next_sum_iv_2[18] ));
    NOR2 inf_abs2_a_0_I_21 (.A(integral[12]), .B(integral[13]), .Y(
        \DWACT_FINC_E[3] ));
    AO1A \preg_RNIUL8B1[16]  (.A(\preg[16]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[16] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I418_Y_0 (.A(sum_0_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I418_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I87_Y (.A(N514), .B(N517), .Y(
        N637));
    AO1 \preg_RNISL4J1[11]  (.A(\preg[11]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[11] ), .Y(
        \un1_next_sum_iv_1[11] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I384_Y_2 (.A(
        ADD_40x40_fast_I384_Y_0), .B(I278_un1_Y), .C(I384_un1_Y), .Y(
        ADD_40x40_fast_I384_Y_2));
    OA1 next_ireg_3_0_ADD_22x22_fast_I29_Y (.A(\i_adj[14]_net_1 ), .B(
        \i_adj[16]_net_1 ), .C(N306), .Y(N334));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I22_P0N (.A(\un1_next_sum[22] ), 
        .B(sum_22), .Y(N538));
    NOR3A inf_abs1_a_2_I_31 (.A(\DWACT_FINC_E[6] ), .B(sr_new[9]), .C(
        sr_new[10]), .Y(N_3));
    OA1 next_ireg_3_0_ADD_22x22_fast_I27_Y (.A(\i_adj[14]_net_1 ), .B(
        \i_adj[16]_net_1 ), .C(N312), .Y(N332));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I223_Y (.A(N700), .B(N708), .Y(
        N782));
    OR2 \ireg_RNIIDF92[25]  (.A(\un1_next_sum_0_iv_1[25] ), .B(
        \ireg_m[25] ), .Y(\un1_next_sum_0_iv[25] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I2_P0N (.A(sum_2_d0), .B(
        \un1_next_sum[0] ), .Y(N478));
    DFN1E1C0 \ireg[6]  (.D(\next_ireg_3[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[6]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I127_un1_Y_0 (.A(N381), .B(N373)
        , .Y(ADD_22x22_fast_I127_un1_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I334_un1_Y (.A(N842), .B(N873), 
        .Y(I334_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I349_un1_Y_0 (.A(N792), .B(
        N776), .Y(ADD_40x40_fast_I349_un1_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I294_un1_Y (.A(N797), .B(N782), 
        .Y(I294_un1_Y));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I23_G0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[23] ), .C(sum_23), .Y(N540));
    DFN1E1C0 \preg[6]  (.D(\p_adj[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[6]_net_1 ));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I36_Y (.A(N293), .B(
        \i_adj[12]_net_1 ), .C(\i_adj[10]_net_1 ), .Y(N341));
    NOR2 inf_abs1_a_2_I_6 (.A(sr_new[0]), .B(sr_new[1]), .Y(N_12));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I1_G0N (.A(\i_adj[1]_net_1 ), 
        .B(\i_adj[3]_net_1 ), .Y(N269));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I318_Y (.A(N727), .B(I250_un1_Y), 
        .C(I318_un1_Y), .Y(N1097));
    AO1 next_ireg_3_0_ADD_22x22_fast_I114_Y (.A(N391), .B(N359), .C(
        N390), .Y(N528));
    AO13 un1_sumreg_0_0_ADD_40x40_fast_I64_Y (.A(\sumreg[26]_net_1 ), 
        .B(N546), .C(\un1_next_sum_1_iv[26] ), .Y(N614));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I457_Y_0 (.A(sum_39), .B(
        \un1_next_sum_1_iv[26] ), .Y(ADD_40x40_fast_I457_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I208_un1_Y (.A(N693), .B(N686), 
        .Y(I208_un1_Y));
    XA1B \sumreg_RNO[34]  (.A(N1031), .B(ADD_40x40_fast_I452_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[34] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I81_Y (.A(N354), .B(N350), .Y(
        N389));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I128_Y (.A(N604), .B(N600), .Y(
        N681));
    DFN1E1C0 \sumreg[29]  (.D(\next_sum[29] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[29]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I99_Y (.A(N496), .B(N499), .Y(
        N649));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I169_Y_0 (.A(\i_adj[11]_net_1 ), 
        .B(\i_adj[9]_net_1 ), .Y(ADD_22x22_fast_I169_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I226_Y (.A(N711), .B(N704), .C(
        N703), .Y(N785));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I442_Y_0 (.A(\sumreg[24]_net_1 )
        , .B(\un1_next_sum[24] ), .Y(ADD_40x40_fast_I442_Y_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I212_Y (.A(N608), .B(N612), .C(
        I212_un1_Y), .Y(N771));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I79_Y (.A(sum_19), .B(
        \un1_next_sum[19] ), .C(N526), .Y(N629));
    AO1 next_ireg_3_0_ADD_22x22_fast_I127_Y_0 (.A(N380), .B(N373), .C(
        N372), .Y(ADD_22x22_fast_I127_Y_0));
    OR3 \ireg_RNI81NK1[25]  (.A(next_sum_1_sqmuxa_2), .B(
        next_sum_1_sqmuxa_1), .C(\un3_next_sum_m[25] ), .Y(
        \un1_next_sum_0_iv_1[25] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I167_Y (.A(N639), .B(N643), .Y(
        N720));
    OR2 \preg_RNIROP64[6]  (.A(\un1_next_sum_iv_2[6] ), .B(
        \un1_next_sum_iv_1[6] ), .Y(\un1_next_sum[6] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I164_Y_0 (.A(\i_adj[4]_net_1 ), 
        .B(\i_adj[6]_net_1 ), .Y(ADD_22x22_fast_I164_Y_0));
    NOR3 inf_abs1_a_2_I_10 (.A(sr_new[0]), .B(sr_new[2]), .C(sr_new[1])
        , .Y(\DWACT_FINC_E[0] ));
    DFN1C0 \state_0[3]  (.D(\state[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_0[3]_net_1 ));
    DFN1E1C0 \ireg[21]  (.D(\next_ireg_3[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[21]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I281_Y (.A(N768), .B(N784), .Y(
        N852));
    XNOR2 inf_abs2_a_0_I_32 (.A(integral[17]), .B(N_16), .Y(
        \inf_abs2_a_0[11] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I430_Y_0 (.A(sum_12), .B(
        \un1_next_sum[12] ), .Y(ADD_40x40_fast_I430_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I217_Y (.A(N702), .B(N694), .Y(
        N776));
    NOR3B \ireg_RNIPI601[6]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[6]_net_1 ), .Y(\un3_next_sum_m[6] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I378_un1_Y (.A(N817), .B(N870), 
        .C(N838), .Y(I378_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I275_Y (.A(N762), .B(N778), .Y(
        N846));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I15_P0N (.A(\un1_next_sum[15] ), 
        .B(sum_15), .Y(N517));
    XA1B \sumreg_RNO[27]  (.A(N1049), .B(ADD_40x40_fast_I445_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[27] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I74_Y (.A(N347), .B(N344), .C(
        N343), .Y(N382));
    DFN1E1C0 \sumreg[19]  (.D(\next_sum[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_19));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I422_Y_0 (.A(sum_4), .B(
        \un1_next_sum[4] ), .Y(ADD_40x40_fast_I422_Y_0));
    DFN1E1C0 \sumreg[8]  (.D(\next_sum[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_8));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I353_un1_Y (.A(
        ADD_40x40_fast_I353_un1_Y_0), .B(N1106), .Y(I353_un1_Y));
    DFN1E1C0 \sumreg[28]  (.D(\next_sum[28] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[28]_net_1 ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I179_Y_0 (.A(\i_adj[21]_net_1 ), 
        .B(\i_adj[19]_net_1 ), .Y(ADD_22x22_fast_I179_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_3 (.A(
        ADD_22x22_fast_I142_un1_Y_0), .B(N421), .C(
        ADD_22x22_fast_I142_Y_2), .Y(ADD_22x22_fast_I142_Y_3));
    XA1B \sumreg_RNO[0]  (.A(N_228), .B(ADD_40x40_fast_I418_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[0] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I256_un1_Y (.A(N741), .B(N734), 
        .Y(I256_un1_Y));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I451_Y_0 (.A(
        \sumreg[33]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I451_Y_0));
    OR2 un1_sumreg_0_0_ADD_m8_i_1 (.A(N_228_1), .B(ADD_m8_i_a4_0_0), 
        .Y(ADD_m8_i_1));
    AO1 \preg_RNILF5Q1[6]  (.A(\preg[6]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[6] ), .Y(
        \un1_next_sum_iv_1[6] ));
    NOR3B \ireg_RNIRK601[8]  (.A(integral[25]), .B(\state[3]_net_1 ), 
        .C(\ireg[8]_net_1 ), .Y(\un3_next_sum_m[8] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I143_Y (.A(N615), .B(N619), .Y(
        N696));
    NOR3B \ireg_RNI78KQ[15]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[15]_net_1 ), .Y(\un3_next_sum_m[15] ));
    DFN1C0 \state_2[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_2[2]_net_1 ));
    DFN1E1C0 \sumreg[18]  (.D(\next_sum[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_18));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I380_Y_1 (.A(N598), .B(N594), .C(
        N683), .Y(ADD_40x40_fast_I380_Y_1));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I61_Y (.A(\sumreg[28]_net_1 ), 
        .B(\sumreg[27]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N611)
        );
    NOR2B next_ireg_3_0_ADD_22x22_fast_I6_G0N (.A(\i_adj[6]_net_1 ), 
        .B(\i_adj[8]_net_1 ), .Y(N284));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I162_Y (.A(
        ADD_22x22_fast_I162_Y_0), .B(N359), .Y(\next_ireg_3[8] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I21_P0N (.A(\un1_next_sum[21] ), 
        .B(sum_21), .Y(N535));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I243_Y (.A(N728), .B(N720), .Y(
        N802));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I127_Y (.A(N603), .B(N599), .Y(
        N680));
    DFN1E1C0 \p_adj[3]  (.D(\inf_abs1_5[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[3]_net_1 ));
    DFN1E1C0 \ireg[10]  (.D(\next_ireg_3[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[10]_net_1 ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I49_Y (.A(\i_adj[3]_net_1 ), .B(
        \i_adj[5]_net_1 ), .C(N279), .Y(N354));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I65_Y (.A(N550), .B(N547), .Y(
        N615));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I47_Y (.A(N279), .B(N282), .Y(
        N352));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I101_Y (.A(N493), .B(N496), .Y(
        N651));
    AND3 inf_abs2_a_0_I_22 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_19));
    AO1 \preg_RNIQJ4J1[10]  (.A(\preg[10]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[10] ), .Y(
        \un1_next_sum_iv_1[10] ));
    OR2 \ireg_RNI3SJQ1[22]  (.A(\un1_next_sum_iv_0[22] ), .B(N_228_1), 
        .Y(\un1_next_sum[22] ));
    DFN1E1C0 \sumreg[1]  (.D(\next_sum[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_1_d0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I449_Y_0 (.A(
        \sumreg[31]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I449_Y_0));
    XA1B \sumreg_RNO[20]  (.A(N1070), .B(ADD_40x40_fast_I438_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[20] ));
    DFN1E1C0 \sumreg_0[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(sum_0_0));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I47_Y (.A(\sumreg[34]_net_1 ), 
        .B(\sumreg[35]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N597)
        );
    XNOR2 inf_abs1_a_2_I_32 (.A(sr_new[11]), .B(N_3), .Y(
        \inf_abs1_a_2[11] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I148_Y (.A(N624), .B(N621), .C(
        N620), .Y(N701));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I165_Y (.A(
        ADD_22x22_fast_I165_Y_0), .B(N531), .Y(\next_ireg_3[11] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I13_G0N (.A(\un1_next_sum[13] )
        , .B(sum_13), .Y(N510_0));
    XA1B \sumreg_RNO[21]  (.A(N1067), .B(ADD_40x40_fast_I439_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[21] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I250_un1_Y (.A(N735), .B(N728), 
        .Y(I250_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I131_Y (.A(N607), .B(N603), .Y(
        N684));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I86_un1_Y (.A(N356), .B(N359), 
        .Y(I86_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I303_Y (.A(N806), .B(N790), .Y(
        N874));
    XNOR2 inf_abs1_a_2_I_20 (.A(sr_new[7]), .B(N_7_0), .Y(
        \inf_abs1_a_2[7] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I438_Y_0 (.A(N_228_1), .B(
        \un1_next_sum_iv_0[20] ), .C(sum_20), .Y(
        ADD_40x40_fast_I438_Y_0));
    DFN1E1C0 \sumreg[25]  (.D(\next_sum[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[25]_net_1 ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I246_Y (.A(I246_un1_Y), .B(N723), 
        .Y(N805));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I151_Y (.A(N623), .B(N627), .Y(
        N704));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I176_Y (.A(N652), .B(N649), .C(
        N648), .Y(N729));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I347_Y (.A(
        ADD_40x40_fast_I347_un1_Y_0), .B(N1088), .C(
        ADD_40x40_fast_I347_Y_0), .Y(N1040));
    DFN1E1C0 \ireg[23]  (.D(\next_ireg_3[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[23]_net_1 ));
    AO1 \preg_RNIUN4J1[12]  (.A(\preg[12]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[12] ), .Y(
        \un1_next_sum_iv_1[12] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I429_Y_0 (.A(
        \un1_next_sum_iv_1[11] ), .B(\un1_next_sum_iv_2[11] ), .C(
        sum_11), .Y(ADD_40x40_fast_I429_Y_0));
    OR2 un1_sumreg_0_0_ADD_m8_i (.A(ADD_m8_i_1), .B(ADD_m8_i_a4_2), .Y(
        N743));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I9_G0N (.A(
        \un1_next_sum_iv_1[9] ), .B(\un1_next_sum_iv_2[9] ), .C(sum_9), 
        .Y(N498));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I142_un1_Y_0 (.A(N373), .B(N365)
        , .C(N396), .Y(ADD_22x22_fast_I142_un1_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I447_Y_0 (.A(
        \sumreg[29]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I447_Y_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I353_Y (.A(I296_un1_Y), .B(N783), 
        .C(I353_un1_Y), .Y(N1058));
    OR2 \ireg_RNI9PUE3[15]  (.A(\un1_next_sum_iv_2[15] ), .B(
        \un1_next_sum_iv_1[15] ), .Y(\un1_next_sum[15] ));
    NOR3B \ireg_RNI8DRU[24]  (.A(integral_1_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[24]_net_1 ), .Y(\un3_next_sum_m[24] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I379_Y_4 (.A(N840), .B(N871), .C(
        ADD_40x40_fast_I379_Y_3), .Y(ADD_40x40_fast_I379_Y_4));
    OR2 next_ireg_3_0_ADD_22x22_fast_I17_P0N (.A(\i_adj[19]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(N318));
    AND3 inf_abs2_a_0_I_60 (.A(integral_i[24]), .B(integral_i[25]), .C(
        integral_i[25]), .Y(\DWACT_FINC_E[15] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I170_Y (.A(N646), .B(N643), .C(
        N642), .Y(N723));
    DFN1E1C0 \sumreg[15]  (.D(\next_sum[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_15));
    DFN1E1C0 \ireg[5]  (.D(\i_adj[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[5]_net_1 ));
    DFN1E1C0 \ireg[25]  (.D(\next_ireg_3[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[25]_net_1 ));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I142_Y_0 (.A(\i_adj[18]_net_1 ), 
        .B(\i_adj[20]_net_1 ), .C(N317), .Y(ADD_22x22_fast_I142_Y_0));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I5_G0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[5] ), .C(sum_5), .Y(N486));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I427_Y_0 (.A(
        \un1_next_sum_iv_1[9] ), .B(\un1_next_sum_iv_2[9] ), .C(sum_9), 
        .Y(ADD_40x40_fast_I427_Y_0));
    DFN1E1C0 \p_adj[9]  (.D(\inf_abs1_5[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[9]_net_1 ));
    XNOR2 inf_abs1_a_2_I_17 (.A(sr_new[6]), .B(N_8_0), .Y(
        \inf_abs1_a_2[6] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I163_Y (.A(
        ADD_22x22_fast_I163_Y_0), .B(N396), .Y(\next_ireg_3[9] ));
    MX2 \i_adj_RNO[14]  (.A(integral[20]), .B(\inf_abs2_a_0[14] ), .S(
        integral_1_0), .Y(\inf_abs2_5[14] ));
    NOR3 \state_RNIRMFQ[6]  (.A(sum_rdy), .B(\state[6]_net_1 ), .C(
        \state[1]_net_1 ), .Y(N_416));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I69_Y (.A(\sumreg[24]_net_1 ), 
        .B(\un1_next_sum[24] ), .C(N541), .Y(N619));
    XA1B \sumreg_RNO[14]  (.A(N1088), .B(ADD_40x40_fast_I432_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[14] ));
    XA1B \sumreg_RNO[35]  (.A(N1029), .B(ADD_40x40_fast_I453_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[35] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I349_Y (.A(
        ADD_40x40_fast_I349_un1_Y_0), .B(N1094), .C(
        ADD_40x40_fast_I349_Y_0), .Y(N1046));
    DFN1C0 \state[4]  (.D(\state[3]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[4]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I147_Y (.A(N619), .B(N623), .Y(
        N700));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I8_G0N (.A(\i_adj[8]_net_1 ), 
        .B(\i_adj[10]_net_1 ), .Y(N290));
    OR2 next_ireg_3_0_ADD_22x22_fast_I9_P0N (.A(\i_adj[9]_net_1 ), .B(
        \i_adj[11]_net_1 ), .Y(N294));
    DFN1E1C0 \sumreg[26]  (.D(\next_sum[26] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[26]_net_1 ));
    OR2 \ireg_RNI7N193[14]  (.A(\un1_next_sum_iv_2[14] ), .B(
        \un1_next_sum_iv_1[14] ), .Y(\un1_next_sum[14] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I441_Y_0 (.A(N_228_1), .B(
        \un1_next_sum_iv_0[23] ), .C(sum_23), .Y(
        ADD_40x40_fast_I441_Y_0));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I179_Y (.A(N490), .B(N487), .C(
        N651), .Y(N732));
    XA1B \sumreg_RNO[7]  (.A(N817), .B(ADD_40x40_fast_I425_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[7] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I11_P0N (.A(
        \un1_next_sum_iv_1[11] ), .B(\un1_next_sum_iv_2[11] ), .C(
        sum_11), .Y(N505));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I267_Y (.A(N754), .B(N770), .Y(
        N838));
    AO1 next_ireg_3_0_ADD_22x22_fast_I128_Y_0 (.A(N382), .B(N375), .C(
        N374), .Y(ADD_22x22_fast_I128_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I90_Y (.A(N507_0), .B(N511), .C(
        N510_0), .Y(N640));
    DFN1E1C0 \ireg[17]  (.D(\next_ireg_3[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[17]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I316_Y (.A(N806), .B(N821), .C(
        N805), .Y(N1091));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I305_Y (.A(N808), .B(N792), .Y(
        N876));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I381_Y (.A(
        ADD_40x40_fast_I381_Y_2), .B(I381_un1_Y), .C(I336_un1_Y), .Y(
        N1027));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I219_Y (.A(N704), .B(N696), .Y(
        N778));
    AO1A \preg_RNISJ8B1[14]  (.A(\preg[14]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[14] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I102_Y (.A(N489), .B(N493), .C(
        N492), .Y(N652));
    NOR2B un1_sumreg_0_0_ADD_m8_i_a4_0_1 (.A(sum_2_d0), .B(
        ADD_m8_i_a4_0_0_0), .Y(ADD_m8_i_a4_0_1));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I70_Y (.A(I70_un1_Y), .B(N540), 
        .Y(N620));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I21_G0N (.A(\un1_next_sum[21] )
        , .B(sum_21), .Y(N534));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I195_Y (.A(
        ADD_40x40_fast_I195_Y_1), .B(N680), .Y(N754));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I421_Y_0 (.A(sum_3), .B(N743), 
        .Y(ADD_40x40_fast_I421_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I318_un1_Y (.A(N810), .B(N743), 
        .Y(I318_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I174_Y (.A(N650), .B(N647), .C(
        N646), .Y(N727));
    DFN1E1C0 \sumreg[16]  (.D(\next_sum[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_16));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I16_G0N (.A(\i_adj[16]_net_1 ), 
        .B(\i_adj[18]_net_1 ), .Y(N314));
    XNOR2 inf_abs2_a_0_I_14 (.A(integral[11]), .B(N_22), .Y(
        \inf_abs2_a_0[5] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I355_Y (.A(N872), .B(N819), .C(
        N871), .Y(N1064));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I132_Y (.A(N608), .B(N604), .Y(
        N685));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I2_G0N (.A(\i_adj[2]_net_1 ), 
        .B(\i_adj[4]_net_1 ), .Y(N272));
    NOR3B \ireg_RNIATL41[7]  (.A(\state[3]_net_1 ), .B(\ireg[7]_net_1 )
        , .C(integral_1_0), .Y(\ireg_m[7] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I152_Y (.A(N628), .B(N625), .C(
        N624), .Y(N705));
    MX2 \p_adj_RNO[8]  (.A(sr_new[8]), .B(\inf_abs1_a_2[8] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[8] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I3_P0N (.A(sum_3), .B(
        \un1_next_sum[0] ), .Y(N481));
    AO1 next_ireg_3_0_ADD_22x22_fast_I76_Y (.A(N349), .B(N346), .C(
        N345), .Y(N384));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I352_un1_Y (.A(
        ADD_40x40_fast_I352_un1_Y_0), .B(N1103), .Y(I352_un1_Y));
    DFN1E1C0 \sumreg[21]  (.D(\next_sum[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(sum_21));
    AO1 next_ireg_3_0_ADD_22x22_fast_I127_Y (.A(
        ADD_22x22_fast_I127_un1_Y_0), .B(N525), .C(
        ADD_22x22_fast_I127_Y_0), .Y(N501));
    XA1 \ireg_RNI8RL41[5]  (.A(integral_1_0), .B(\ireg[5]_net_1 ), .C(
        \state[3]_net_1 ), .Y(\un1_next_sum_iv_0[5] ));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I143_un1_Y (.A(N423), .B(N407), 
        .C(N359), .Y(I143_un1_Y));
    MX2 \p_adj_RNO[7]  (.A(sr_new[7]), .B(\inf_abs1_a_2[7] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[7] ));
    XA1 \ireg_RNI68LQ[23]  (.A(integral_0_0), .B(\ireg[23]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[23] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I84_Y (.A(N516), .B(N520), .C(
        N519), .Y(N634));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I42_Y (.A(N284), .B(
        \i_adj[9]_net_1 ), .C(\i_adj[7]_net_1 ), .Y(N347));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I222_Y (.A(N707), .B(N700), .C(
        N699), .Y(N781));
    XA1B \sumreg_RNO[36]  (.A(N1027), .B(ADD_40x40_fast_I454_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[36] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I1_P0N (.A(sum_1_d0), .B(
        \un1_next_sum[0] ), .Y(N475));
    OA1 next_ireg_3_0_ADD_22x22_fast_I31_Y (.A(\i_adj[12]_net_1 ), .B(
        \i_adj[14]_net_1 ), .C(N306), .Y(N336));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I70_un1_Y (.A(sum_22), .B(
        \un1_next_sum[22] ), .C(N541), .Y(I70_un1_Y));
    OR2 \preg_RNISE1P3[12]  (.A(\un1_next_sum_iv_2[12] ), .B(
        \un1_next_sum_iv_1[12] ), .Y(\un1_next_sum[12] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I129_Y (.A(
        ADD_22x22_fast_I129_un1_Y_0), .B(N531), .C(
        ADD_22x22_fast_I129_Y_0), .Y(N507));
    OR3 next_ireg_3_0_ADD_22x22_fast_I143_Y (.A(I143_un1_Y), .B(
        ADD_22x22_fast_I143_Y_2), .C(I122_un1_Y), .Y(N494));
    DFN1E1C0 \p_adj[1]  (.D(\inf_abs1_5[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[1]_net_1 ));
    NOR3A inf_abs1_a_2_I_27 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .C(
        sr_new[9]), .Y(N_4));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I186_Y (.A(N662), .B(N659), .C(
        N658), .Y(N739));
    OR2 \state_RNIFG0J1[3]  (.A(N_228_1), .B(next_sum_0_sqmuxa), .Y(
        \un1_next_sum[0] ));
    NOR2 inf_abs2_a_0_I_15 (.A(integral[9]), .B(integral[10]), .Y(
        \DWACT_FINC_E[1] ));
    AX1D un1_sumreg_0_0_ADD_40x40_fast_I434_Y_0 (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(ADD_40x40_fast_I434_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I227_Y (.A(N704), .B(N712), .Y(
        N786));
    DFN1E1C0 \p_adj[7]  (.D(\inf_abs1_5[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[7]_net_1 ));
    NOR2B \preg_RNIVKAK[18]  (.A(\preg[18]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[18] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I299_Y (.A(N802), .B(N786), .Y(
        N870));
    DFN1E1C0 \sumreg[11]  (.D(\next_sum[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_11));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I433_Y_0 (.A(sum_15), .B(
        \un1_next_sum[15] ), .Y(ADD_40x40_fast_I433_Y_0));
    XA1B \sumreg_RNO[33]  (.A(N1033), .B(ADD_40x40_fast_I451_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[33] ));
    DFN1E1C0 \ireg[19]  (.D(\next_ireg_3[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[19]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I320_un1_Y (.A(N814), .B(N666), 
        .Y(I320_un1_Y));
    MX2 \i_adj_RNO[10]  (.A(integral[16]), .B(\inf_abs2_a_0[10] ), .S(
        integral_1_0), .Y(\inf_abs2_5[10] ));
    XNOR2 inf_abs2_a_0_I_40 (.A(integral[20]), .B(N_13), .Y(
        \inf_abs2_a_0[14] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I385_Y_0 (.A(N685), .B(
        I208_un1_Y), .Y(ADD_40x40_fast_I385_Y_0));
    AND3 inf_abs2_a_0_I_54 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E[9] ), .C(\DWACT_FINC_E[12] ), .Y(
        \DWACT_FINC_E[13] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I180_Y (.A(N656), .B(N653), .C(
        N652), .Y(N733));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I167_Y (.A(\i_adj[7]_net_1 ), .B(
        \i_adj[9]_net_1 ), .C(N525), .Y(\next_ireg_3[13] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I57_Y (.A(\sumreg[29]_net_1 ), 
        .B(\sumreg[30]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N607)
        );
    DFN1C0 \state[1]  (.D(\state_RNIGPKC[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state[1]_net_1 ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I382_Y (.A(
        ADD_40x40_fast_I382_Y_1), .B(I382_un1_Y), .C(I338_un1_Y), .Y(
        N1029));
    MX2 \p_adj_RNO[10]  (.A(sr_new[10]), .B(\inf_abs1_a_2[10] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[10] ));
    DFN1E1C0 \ireg[22]  (.D(\next_ireg_3[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[22]_net_1 ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I20_P0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[20] ), .C(sum_20), .Y(N532));
    AX1D next_ireg_3_0_ADD_22x22_fast_I169_Y (.A(N424), .B(I133_un1_Y), 
        .C(ADD_22x22_fast_I169_Y_0), .Y(\next_ireg_3[15] ));
    OR2A un1_sumreg_0_0_ADD_40x40_fast_I37_P0N (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[37]_net_1 ), .Y(N583));
    NOR3B inf_abs2_a_0_I_16 (.A(\DWACT_FINC_E[1] ), .B(
        \DWACT_FINC_E_0[0] ), .C(integral[11]), .Y(N_21));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I278_un1_Y (.A(N692), .B(N684), 
        .C(N781), .Y(I278_un1_Y));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_1 (.A(N326), .B(N329), .C(
        ADD_22x22_fast_I142_Y_0), .Y(ADD_22x22_fast_I142_Y_1));
    NOR3B inf_abs2_a_0_I_55 (.A(\DWACT_FINC_E[13] ), .B(
        \DWACT_FINC_E[28] ), .C(integral[24]), .Y(N_8));
    DFN1E1C0 \preg[13]  (.D(\p_adj[7]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[13]_net_1 ));
    AO1 \preg_RNIRL5Q1[9]  (.A(\preg[9]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[9] ), .Y(
        \un1_next_sum_iv_1[9] ));
    DFN1E1C0 \i_adj[6]  (.D(\inf_abs2_5[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[6]_net_1 ));
    DFN1E1C0 \i_adj[4]  (.D(\inf_abs2_5[4] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[4]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I63_Y (.A(N336), .B(N332), .Y(
        N371));
    NOR2B un1_sumreg_0_0_ADD_m8_i_a4_0 (.A(ADD_m8_i_a4_0_1), .B(N_232), 
        .Y(ADD_m8_i_a4_0_0));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I230_Y (.A(I230_un1_Y), .B(N707), 
        .Y(N789));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I81_Y (.A(sum_17), .B(
        \un1_next_sum[17] ), .C(N526), .Y(N631));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I379_Y_2 (.A(N596), .B(
        ADD_40x40_fast_I379_Y_0), .C(N681), .Y(ADD_40x40_fast_I379_Y_2)
        );
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I230_un1_Y (.A(N715), .B(N708), 
        .Y(I230_un1_Y));
    MX2 \i_adj_RNO[18]  (.A(integral[24]), .B(\inf_abs2_a_0[18] ), .S(
        integral[25]), .Y(\inf_abs2_5[18] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I456_Y_0 (.A(
        \sumreg[38]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I456_Y_0));
    NOR2A inf_abs1_a_2_I_11 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .Y(
        N_10));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I348_Y (.A(I286_un1_Y), .B(N773), 
        .C(I348_un1_Y), .Y(N1043));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I165_Y (.A(N637), .B(N641), .Y(
        N718));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I381_Y_1 (.A(N600), .B(N596), .C(
        N685), .Y(ADD_40x40_fast_I381_Y_1));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I92_Y (.A(N504_0), .B(sum_12), 
        .C(\un1_next_sum[12] ), .Y(N642));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I348_un1_Y (.A(N774), .B(N790), 
        .C(N1091), .Y(I348_un1_Y));
    DFN1E1C0 \i_adj[9]  (.D(\inf_abs2_5[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[9]_net_1 ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I182_un1_Y (.A(N490), .B(N487), 
        .C(N658), .Y(I182_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I85_Y (.A(N517), .B(N520), .Y(
        N635));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I11_G0N (.A(
        \un1_next_sum_iv_1[11] ), .B(\un1_next_sum_iv_2[11] ), .C(
        sum_11), .Y(N504_0));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I201_Y (.A(N597), .B(N601), .C(
        N686), .Y(N760));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I72_Y (.A(N534), .B(sum_22), .C(
        \un1_next_sum[22] ), .Y(N622));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I0_S (.A(\i_adj[0]_net_1 ), .B(
        \i_adj[2]_net_1 ), .Y(\next_ireg_3[6] ));
    NOR3C next_ireg_3_0_ADD_22x22_fast_I120_un1_Y (.A(N373), .B(N365), 
        .C(N420), .Y(I120_un1_Y));
    DFN1E1C0 \i_adj[3]  (.D(\inf_abs2_5[3] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[3]_net_1 ));
    XA1B \sumreg_RNO[15]  (.A(N1085), .B(ADD_40x40_fast_I433_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[15] ));
    NOR3B \ireg_RNI6AQU[13]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[13]_net_1 ), .C(integral_1_0), .Y(\ireg_m[13] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I242_Y (.A(I242_un1_Y), .B(N719), 
        .Y(N801));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y_1 (.A(N371), .B(N378), .C(
        ADD_22x22_fast_I126_Y_0), .Y(ADD_22x22_fast_I126_Y_1));
    OA1 next_ireg_3_0_ADD_22x22_fast_I51_Y (.A(\i_adj[3]_net_1 ), .B(
        \i_adj[5]_net_1 ), .C(N273), .Y(N356));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I178_Y (.A(\i_adj[18]_net_1 ), 
        .B(\i_adj[20]_net_1 ), .C(N494), .Y(\next_ireg_3[24] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I231_Y (.A(N708), .B(N716), .Y(
        N790));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I184_Y (.A(I184_un1_Y), .B(N656), 
        .Y(N737));
    XNOR2 inf_abs2_a_0_I_56 (.A(integral[25]), .B(N_8), .Y(
        \inf_abs2_a_0[19] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I87_Y (.A(I87_un1_Y), .B(N357), 
        .Y(N396));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I251_Y (.A(N736), .B(N728), .Y(
        N810));
    DFN1E1C0 \sumreg[34]  (.D(\next_sum[34] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[34]_net_1 ));
    AO1A \ireg_RNI81002[16]  (.A(\ireg[16]_net_1 ), .B(
        next_sum_0_sqmuxa), .C(\un1_next_sum_iv_0[16] ), .Y(
        \un1_next_sum_iv_2[16] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I340_un1_Y (.A(N795), .B(
        I308_un1_Y), .C(N848), .Y(I340_un1_Y));
    AO1 \ireg_RNI3Q191[14]  (.A(\ireg[14]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[14] ), .Y(
        \un1_next_sum_iv_1[14] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I247_Y (.A(N732), .B(N724), .Y(
        N806));
    DFN1C0 \state_0[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_0[2]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I60_Y (.A(\sumreg[27]_net_1 ), 
        .B(\sumreg[28]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N610)
        );
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I385_un1_Y (.A(N884), .B(
        \un1_next_sum[0] ), .C(N852), .Y(I385_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I173_Y (.A(N649), .B(N645), .Y(
        N726));
    OR2 next_ireg_3_0_ADD_22x22_fast_I6_P0N (.A(\i_adj[6]_net_1 ), .B(
        \i_adj[8]_net_1 ), .Y(N285));
    DFN1E1C0 \ireg[7]  (.D(\next_ireg_3[7] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[7]_net_1 ));
    XA1B \sumreg_RNO[28]  (.A(N1046), .B(ADD_40x40_fast_I446_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[28] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I380_un1_Y (.A(N821), .B(N874), 
        .C(N842), .Y(I380_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I238_Y (.A(N723), .B(N716), .C(
        N715), .Y(N797));
    XA1B \sumreg_RNO[3]  (.A(\un1_next_sum[0] ), .B(
        ADD_40x40_fast_I421_Y_0), .C(\state_2[2]_net_1 ), .Y(
        \next_sum[3] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I269_Y (.A(N756), .B(N772), .Y(
        N840));
    DFN1E1C0 \preg[7]  (.D(\p_adj[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[7]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I44_Y (.A(\sumreg[36]_net_1 ), 
        .B(\sumreg[35]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N594)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I258_Y (.A(N736), .B(N743), .C(
        N735), .Y(N817));
    DFN1E1C0 \ireg[16]  (.D(\next_ireg_3[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[16]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I273_Y (.A(N760), .B(N776), .Y(
        N844));
    AND2 un1_sumreg_0_0_ADD_40x40_fast_I195_Y_0 (.A(N583), .B(N586), 
        .Y(ADD_40x40_fast_I195_Y_0));
    XA1B \sumreg_RNO[32]  (.A(N1035), .B(ADD_40x40_fast_I450_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[32] ));
    DFN1E1C0 \preg[10]  (.D(\p_adj[4]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[10]_net_1 ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I163_Y_0 (.A(\i_adj[3]_net_1 ), 
        .B(\i_adj[5]_net_1 ), .Y(ADD_22x22_fast_I163_Y_0));
    DFN1E1C0 \preg[18]  (.D(\p_adj[12]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[18]_net_1 ));
    AND2 \un1_next_sum_iv_0_RNO_0[19]  (.A(next_sum_1_sqmuxa), .B(
        \ireg[19]_net_1 ), .Y(\ireg_m[19] ));
    NOR3 inf_abs2_a_0_I_18 (.A(integral[10]), .B(integral[9]), .C(
        integral[11]), .Y(\DWACT_FINC_E[2] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I6_P0N (.A(\un1_next_sum[6] ), 
        .B(sum_6), .Y(N490));
    XA1B \sumreg_RNO[8]  (.A(N1106), .B(ADD_40x40_fast_I426_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[8] ));
    NOR2B \preg_RNISHAK[15]  (.A(\preg[15]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[15] ));
    OA1 next_ireg_3_0_ADD_22x22_fast_I23_Y (.A(\i_adj[18]_net_1 ), .B(
        \i_adj[16]_net_1 ), .C(N318), .Y(N328));
    AND2 \un1_next_sum_iv_0_RNO_0[21]  (.A(next_sum_1_sqmuxa), .B(
        \ireg[21]_net_1 ), .Y(\ireg_m[21] ));
    AO1A \preg_RNIGPDC1[9]  (.A(\preg[9]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[9] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I178_Y (.A(N654), .B(N651), .C(
        N650), .Y(N731));
    NOR2B inf_abs2_a_0_I_34 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .Y(N_15));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I98_Y (.A(N495), .B(N499), .C(
        N498), .Y(N648));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I7_P0N (.A(\un1_next_sum[7] ), 
        .B(sum_7), .Y(N493));
    NOR2 inf_abs2_a_0_I_47 (.A(integral[21]), .B(integral[22]), .Y(
        \DWACT_FINC_E[11] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I89_Y (.A(N514), .B(N511), .Y(
        N639));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I10_P0N (.A(\un1_next_sum[10] ), 
        .B(sum_10), .Y(N502));
    NOR2 inf_abs1_a_2_I_21 (.A(sr_new[6]), .B(sr_new[7]), .Y(
        \DWACT_FINC_E_0[3] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I5_G0N (.A(\i_adj[7]_net_1 ), 
        .B(\i_adj[5]_net_1 ), .Y(N281));
    AX1D next_ireg_3_0_ADD_22x22_fast_I176_Y (.A(I126_un1_Y), .B(
        ADD_22x22_fast_I126_Y_1), .C(ADD_22x22_fast_I176_Y_0), .Y(
        \next_ireg_3[22] ));
    NOR3 inf_abs2_a_0_I_8 (.A(integral[7]), .B(integral[6]), .C(
        integral[8]), .Y(N_24));
    XA1B \sumreg_RNO[16]  (.A(N1082), .B(ADD_40x40_fast_I434_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[16] ));
    NOR3B inf_abs2_a_0_I_19 (.A(\DWACT_FINC_E[2] ), .B(
        \DWACT_FINC_E_0[0] ), .C(integral[12]), .Y(N_20));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I78_Y (.A(N525_0), .B(sum_19), 
        .C(\un1_next_sum[19] ), .Y(N628));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I132_un1_Y (.A(N423), .B(N359), 
        .Y(I132_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I0_CO1 (.A(\i_adj[0]_net_1 ), 
        .B(\i_adj[2]_net_1 ), .Y(N266));
    OR2A un1_sumreg_0_0_ADD_40x40_fast_I26_P0N (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[26]_net_1 ), .Y(N550));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I65_Y (.A(N334), .B(N338), .Y(
        N373));
    AO1 \preg_RNI0Q4J1[13]  (.A(\preg[13]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[13] ), .Y(
        \un1_next_sum_iv_1[13] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I229_Y (.A(N714), .B(N706), .Y(
        N788));
    XA1B \sumreg_RNO[13]  (.A(N1091), .B(ADD_40x40_fast_I431_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[13] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I112_un1_Y (.A(N387), .B(N394), 
        .Y(I112_un1_Y));
    XNOR2 inf_abs2_a_0_I_7 (.A(integral[8]), .B(N_25), .Y(
        \inf_abs2_a_0[2] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I133_un1_Y (.A(N425), .B(N266), 
        .Y(I133_un1_Y));
    XNOR2 inf_abs2_a_0_I_35 (.A(integral[18]), .B(N_15), .Y(
        \inf_abs2_a_0[12] ));
    OR3 \preg_RNI8BKC2[7]  (.A(\un24_next_sum_m[7] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[7] ), .Y(
        \un1_next_sum_iv_2[7] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I1_P0N (.A(\i_adj[1]_net_1 ), .B(
        \i_adj[3]_net_1 ), .Y(N270));
    XOR2 inf_abs2_a_0_I_5 (.A(integral[6]), .B(integral[7]), .Y(
        \inf_abs2_a_0[1] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I107_Y (.A(N389), .B(N381), .Y(
        N421));
    AND3 inf_abs2_a_0_I_61 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[15] ), .Y(N_6));
    AND3 inf_abs2_a_0_I_58 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[14] ), .Y(N_7));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I111_Y (.A(N481), .B(N478), .Y(
        N661));
    XA1B \sumreg_RNO[19]  (.A(N1073), .B(ADD_40x40_fast_I437_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[19] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I68_Y (.A(N341), .B(N338), .C(
        N337), .Y(N376));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I16_G0N (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(N519));
    XNOR2 inf_abs1_a_2_I_12 (.A(sr_new[4]), .B(N_10), .Y(
        \inf_abs1_a_2[4] ));
    AO1 \preg_RNIPJ5Q1[8]  (.A(\preg[8]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[8] ), .Y(
        \un1_next_sum_iv_1[8] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I446_Y_0 (.A(
        \sumreg[28]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I446_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I109_Y (.A(N391), .B(N383), .Y(
        N423));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I93_Y (.A(sum_12), .B(
        \un1_next_sum[12] ), .C(N505), .Y(N643));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I212_un1_Y (.A(N697), .B(N690), 
        .Y(I212_un1_Y));
    DFN1E1C0 \p_adj[12]  (.D(\inf_abs1_5[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[12]_net_1 ));
    DFN1E1C0 \p_adj[2]  (.D(\inf_abs1_5[2] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[2]_net_1 ));
    MX2 \i_adj_RNO[9]  (.A(integral[15]), .B(\inf_abs2_a_0[9] ), .S(
        integral_0_0), .Y(\inf_abs2_5[9] ));
    DFN1E1C0 \ireg[18]  (.D(\next_ireg_3[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[18]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_1 (.A(N328), .B(N331), .C(
        ADD_22x22_fast_I143_Y_0), .Y(ADD_22x22_fast_I143_Y_1));
    NOR3A inf_abs2_a_0_I_13 (.A(\DWACT_FINC_E_0[0] ), .B(integral[9]), 
        .C(integral[10]), .Y(N_22));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I313_Y (.A(N816), .B(N800), .Y(
        N884));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I73_Y (.A(N535), .B(N538), .Y(
        N623));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I45_Y (.A(\sumreg[35]_net_1 ), 
        .B(\sumreg[36]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N595)
        );
    DFN1E1C0 \ireg[9]  (.D(\next_ireg_3[9] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[9]_net_1 ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I382_Y_0 (.A(N598), .B(N602), .C(
        N687), .Y(ADD_40x40_fast_I382_Y_0));
    DFN1E1C0 \preg[14]  (.D(\p_adj[8]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[14]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I96_Y (.A(N498), .B(N502), .C(
        N501_0), .Y(N646));
    XNOR2 inf_abs2_a_0_I_59 (.A(integral[25]), .B(N_7), .Y(
        \inf_abs2_a_0[20] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I142_Y_2 (.A(N365), .B(N372), .C(
        ADD_22x22_fast_I142_Y_1), .Y(ADD_22x22_fast_I142_Y_2));
    AND3 inf_abs2_a_0_I_24 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E_0[4] ));
    DFN1E1C0 \preg[9]  (.D(\p_adj[3]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[9]_net_1 ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I426_Y_0 (.A(sum_8), .B(
        \un1_next_sum[8] ), .Y(ADD_40x40_fast_I426_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I379_Y (.A(
        ADD_40x40_fast_I379_un1_Y_0), .B(N819), .C(
        ADD_40x40_fast_I379_Y_4), .Y(N1023));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I76_Y (.A(N528_0), .B(N532), .C(
        N531_0), .Y(N626));
    DFN1P0 \state[0]  (.D(\state_ns[0] ), .CLK(clk_c), .PRE(n_rst_c), 
        .Q(sum_rdy));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I205_Y (.A(N682), .B(N690), .Y(
        N764));
    NOR2B inf_abs1_a_2_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_2));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I177_Y (.A(N653), .B(N649), .Y(
        N730));
    NOR3B inf_abs2_a_0_I_36 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .C(integral[18]), .Y(N_14));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I8_G0N (.A(\un1_next_sum[8] ), 
        .B(sum_8), .Y(N495));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I140_un1_Y (.A(N616), .B(N613), 
        .Y(I140_un1_Y));
    XA1B \sumreg_RNO[6]  (.A(N819), .B(ADD_40x40_fast_I424_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[6] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I71_Y (.A(N340), .B(N344), .Y(
        N379));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I145_Y (.A(N617), .B(N621), .Y(
        N698));
    AO1A \state_RNO[0]  (.A(sum_enable), .B(sum_rdy), .C(
        \state[5]_net_1 ), .Y(\state_ns[0] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I62_Y (.A(\sumreg[26]_net_1 ), 
        .B(\sumreg[27]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N612)
        );
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I380_Y (.A(I380_un1_Y), .B(
        ADD_40x40_fast_I380_Y_2), .C(I334_un1_Y), .Y(N1025));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I235_Y (.A(N720), .B(N712), .Y(
        N794));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I191_Y (.A(N472), .B(
        \un1_next_sum[0] ), .C(N664), .Y(N745));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I455_Y_0 (.A(
        \sumreg[37]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I455_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I255_Y (.A(N740), .B(N732), .Y(
        N814));
    AO1 next_ireg_3_0_ADD_22x22_fast_I82_Y (.A(N355), .B(N352), .C(
        N351), .Y(N390));
    NOR2A inf_abs2_a_0_I_25 (.A(\DWACT_FINC_E_0[4] ), .B(integral[14]), 
        .Y(N_18));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I183_Y (.A(N490), .B(N487), .C(
        N659), .Y(N736));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I254_un1_Y (.A(N739), .B(N732), 
        .Y(I254_un1_Y));
    DFN1E1C0 \ireg[8]  (.D(\next_ireg_3[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[8]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I302_un1_Y (.A(N805), .B(N790), 
        .Y(I302_un1_Y));
    OA1 next_ireg_3_0_ADD_22x22_fast_I25_Y (.A(\i_adj[18]_net_1 ), .B(
        \i_adj[16]_net_1 ), .C(N312), .Y(N330));
    OA1 next_ireg_3_0_ADD_22x22_fast_I43_Y (.A(\i_adj[9]_net_1 ), .B(
        \i_adj[7]_net_1 ), .C(N285), .Y(N348));
    XNOR2 inf_abs1_a_2_I_35 (.A(sr_new[12]), .B(N_2), .Y(
        \inf_abs1_a_2[12] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I199_Y_0 (.A(N595), .B(N599), 
        .Y(ADD_40x40_fast_I199_Y_0));
    DFN1E1C0 \preg[8]  (.D(\p_adj[2]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\preg[8]_net_1 ));
    XNOR2 inf_abs2_a_0_I_53 (.A(integral[24]), .B(N_9), .Y(
        \inf_abs2_a_0[18] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I64_Y (.A(N337), .B(N334), .C(
        N333), .Y(N372));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I301_Y (.A(N804), .B(N788), .Y(
        N872));
    DFN1E1C0 \i_adj[14]  (.D(\inf_abs2_5[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[14]_net_1 ));
    DFN1E1C0 \sumreg[32]  (.D(\next_sum[32] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[32]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I346_Y (.A(
        ADD_40x40_fast_I346_un1_Y_0), .B(N1085), .C(
        ADD_40x40_fast_I346_Y_0), .Y(N1037));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I28_Y (.A(N305), .B(
        \i_adj[14]_net_1 ), .C(\i_adj[16]_net_1 ), .Y(N333));
    NOR2A un1_sumreg_0_0_ADD_40x40_fast_I25_G0N (.A(\sumreg[25]_net_1 )
        , .B(\un1_next_sum_0_iv[25] ), .Y(N546));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I249_Y (.A(N734), .B(N726), .Y(
        N808));
    AO1A \ireg_RNIA3002[17]  (.A(\ireg[17]_net_1 ), .B(
        next_sum_0_sqmuxa), .C(\un1_next_sum_iv_0[17] ), .Y(
        \un1_next_sum_iv_2[17] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I351_Y (.A(I292_un1_Y), .B(N779), 
        .C(I351_un1_Y), .Y(N1052));
    MX2 \i_adj_RNO[6]  (.A(integral[12]), .B(\inf_abs2_a_0[6] ), .S(
        integral_0_0), .Y(\inf_abs2_5[6] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I188_Y (.A(N664), .B(N661), .C(
        N660), .Y(N741));
    AND3 inf_abs1_a_2_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(N_6_0));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I16_P0N (.A(
        \un1_next_sum_iv_1[16] ), .B(\un1_next_sum_iv_2[16] ), .C(
        sum_16), .Y(N520));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I49_Y (.A(\sumreg[34]_net_1 ), 
        .B(\sumreg[33]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N599)
        );
    XNOR2 inf_abs2_a_0_I_26 (.A(integral[15]), .B(N_18), .Y(
        \inf_abs2_a_0[9] ));
    XA1B \sumreg_RNO[12]  (.A(N1094), .B(ADD_40x40_fast_I430_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[12] ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I54_Y (.A(\sumreg[30]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N604)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I315_Y (.A(N804), .B(N819), .C(
        N803), .Y(N1088));
    NOR3B \preg_RNIELFL[8]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[8]_net_1 ), .Y(\un24_next_sum_m[8] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I112_Y (.A(sum_1_d0), .B(
        sum_2_d0), .C(\un1_next_sum[0] ), .Y(N662));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I177_Y_0 (.A(\i_adj[19]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(ADD_22x22_fast_I177_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I106_Y (.A(N483), .B(N487), .C(
        N486), .Y(N656));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I7_G0N (.A(\un1_next_sum[7] ), 
        .B(sum_7), .Y(N492));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I242_un1_Y (.A(N727), .B(N720), 
        .Y(I242_un1_Y));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I164_Y (.A(
        ADD_22x22_fast_I164_Y_0), .B(N394), .Y(\next_ireg_3[10] ));
    XNOR2 inf_abs2_a_0_I_62 (.A(integral[25]), .B(N_6), .Y(
        \inf_abs2_a_0[21] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I419_Y_0 (.A(sum_1_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I419_Y_0));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I68_Y (.A(N540), .B(
        \sumreg[24]_net_1 ), .C(\un1_next_sum[24] ), .Y(N618));
    NOR2 inf_abs2_a_0_I_38 (.A(integral[18]), .B(integral[19]), .Y(
        \DWACT_FINC_E[8] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I380_Y_2 (.A(N758), .B(N773), .C(
        ADD_40x40_fast_I380_Y_1), .Y(ADD_40x40_fast_I380_Y_2));
    NOR3 inf_abs2_a_0_I_41 (.A(integral[19]), .B(integral[18]), .C(
        integral[20]), .Y(\DWACT_FINC_E[9] ));
    MX2 \p_adj_RNO[9]  (.A(sr_new[9]), .B(\inf_abs1_a_2[9] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[9] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I162_Y_0 (.A(\i_adj[2]_net_1 ), 
        .B(\i_adj[4]_net_1 ), .Y(ADD_22x22_fast_I162_Y_0));
    NOR2A \ireg_RNIACOK_0[25]  (.A(next_sum_1_sqmuxa), .B(
        \ireg[25]_net_1 ), .Y(\un3_next_sum_m[25] ));
    DFN1E1C0 \sumreg[33]  (.D(\next_sum[33] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[33]_net_1 ));
    XA1B \sumreg_RNO[2]  (.A(N745), .B(ADD_40x40_fast_I420_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[2] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I156_Y (.A(N632), .B(N629), .C(
        N628), .Y(N709));
    NOR3B \preg_RNIDKFL[7]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[7]_net_1 ), .Y(\un24_next_sum_m[7] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I352_un1_Y_0 (.A(N798), .B(
        N782), .Y(ADD_40x40_fast_I352_un1_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I100_Y (.A(N492), .B(N496), .C(
        N495), .Y(N650));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I165_Y_0 (.A(\i_adj[5]_net_1 ), 
        .B(\i_adj[7]_net_1 ), .Y(ADD_22x22_fast_I165_Y_0));
    DFN1E1C0 \i_adj[12]  (.D(\inf_abs2_5[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[12]_net_1 ));
    NOR2B \i_adj_RNO[19]  (.A(\inf_abs2_a_0[19] ), .B(integral[25]), 
        .Y(\inf_abs2_5[19] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I359_un1_Y (.A(N880), .B(N745), 
        .Y(I359_un1_Y));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I39_Y (.A(N291), .B(N294), .Y(
        N344));
    AO1 next_ireg_3_0_ADD_22x22_fast_I126_Y_0 (.A(N335), .B(N332), .C(
        N331), .Y(ADD_22x22_fast_I126_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I14_G0N (.A(\i_adj[16]_net_1 ), 
        .B(\i_adj[14]_net_1 ), .Y(N308));
    AO1A \ireg_RNI4TVV1[14]  (.A(\ireg[14]_net_1 ), .B(
        next_sum_0_sqmuxa), .C(\un1_next_sum_iv_0[14] ), .Y(
        \un1_next_sum_iv_2[14] ));
    DFN1E1C0 \sumreg[30]  (.D(\next_sum[30] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[30]_net_1 ));
    AND3 inf_abs2_a_0_I_39 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E_0[7] ), .C(\DWACT_FINC_E[8] ), .Y(N_13));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I24_Y (.A(N311), .B(
        \i_adj[18]_net_1 ), .C(\i_adj[16]_net_1 ), .Y(N329));
    OA1 next_ireg_3_0_ADD_22x22_fast_I37_Y (.A(\i_adj[12]_net_1 ), .B(
        \i_adj[10]_net_1 ), .C(N294), .Y(N342));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I302_Y (.A(I302_un1_Y), .B(N789), 
        .Y(N873));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I292_un1_Y (.A(N706), .B(N698), 
        .C(N795), .Y(I292_un1_Y));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I130_Y (.A(N606), .B(N602), .Y(
        N683));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I80_Y (.A(N522), .B(N526), .C(
        N525_0), .Y(N630));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I346_un1_Y_0 (.A(N786), .B(
        N770), .Y(ADD_40x40_fast_I346_un1_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I0_G0N (.A(N_228), .B(sum_0_d0)
        , .Y(N471));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I150_Y (.A(I150_un1_Y), .B(N622), 
        .Y(N703));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I161_Y (.A(N637), .B(N633), .Y(
        N714));
    AO1 next_ireg_3_0_ADD_22x22_fast_I40_Y (.A(N287), .B(N291), .C(
        N290), .Y(N345));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I346_Y_0 (.A(N785), .B(N770), .C(
        N769), .Y(ADD_40x40_fast_I346_Y_0));
    OA1A un1_sumreg_0_0_ADD_40x40_fast_I63_Y (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[27]_net_1 ), .C(N550), .Y(
        N613));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I187_Y (.A(N475), .B(N478), .C(
        N659), .Y(N740));
    XA1B \sumreg_RNO[4]  (.A(N823), .B(ADD_40x40_fast_I422_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[4] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I352_Y (.A(I294_un1_Y), .B(N781), 
        .C(I352_un1_Y), .Y(N1055));
    XA1B \sumreg_RNO[5]  (.A(N821), .B(ADD_40x40_fast_I423_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[5] ));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I378_Y (.A(
        ADD_40x40_fast_I378_Y_3), .B(I378_un1_Y), .C(I330_un1_Y), .Y(
        N1021));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I45_Y (.A(N285), .B(N282), .Y(
        N350));
    AX1D next_ireg_3_0_ADD_22x22_fast_I171_Y (.A(N420), .B(I131_un1_Y), 
        .C(ADD_22x22_fast_I171_Y_0), .Y(\next_ireg_3[17] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I432_Y_0 (.A(sum_14), .B(
        \un1_next_sum[14] ), .Y(ADD_40x40_fast_I432_Y_0));
    DFN1E1C0 \sumreg[37]  (.D(\next_sum[37] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[37]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I17_G0N (.A(\i_adj[19]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(N317));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I51_Y (.A(\sumreg[32]_net_1 ), 
        .B(\sumreg[33]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N601)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I383_Y_1 (.A(N764), .B(N779), .C(
        ADD_40x40_fast_I383_Y_0), .Y(ADD_40x40_fast_I383_Y_1));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I23_P0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[23] ), .C(sum_23), .Y(N541));
    AO1 next_ireg_3_0_ADD_22x22_fast_I143_Y_2 (.A(N367), .B(N374), .C(
        ADD_22x22_fast_I143_Y_1), .Y(ADD_22x22_fast_I143_Y_2));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I66_Y (.A(I66_un1_Y), .B(N546), 
        .Y(N616));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I445_Y_0 (.A(
        \sumreg[27]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I445_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I298_un1_Y (.A(N801), .B(N786), 
        .Y(I298_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I109_Y (.A(N481), .B(N484), .Y(
        N659));
    XNOR2 inf_abs2_a_0_I_28 (.A(integral[16]), .B(N_17), .Y(
        \inf_abs2_a_0[10] ));
    NOR3 inf_abs2_a_0_I_33 (.A(integral[16]), .B(integral[15]), .C(
        integral[17]), .Y(\DWACT_FINC_E_0[7] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I55_Y (.A(\sumreg[30]_net_1 ), 
        .B(\sumreg[31]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N605)
        );
    DFN1C0 \state_1[2]  (.D(\state_0[1]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\state_1[2]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I48_Y (.A(N275), .B(N279), .C(
        N278), .Y(N353));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I3_G0N (.A(sum_3), .B(
        \un1_next_sum[0] ), .Y(N480));
    NOR3B \ireg_RNI9SL41[6]  (.A(\state[3]_net_1 ), .B(\ireg[6]_net_1 )
        , .C(integral_1_0), .Y(\ireg_m[6] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I344_un1_Y (.A(N799), .B(
        I312_un1_Y), .C(N852), .Y(I344_un1_Y));
    MX2 \i_adj_RNO[4]  (.A(integral[10]), .B(\inf_abs2_a_0[4] ), .S(
        integral_0_0), .Y(\inf_abs2_5[4] ));
    OR3 \ireg_RNI0PS52[13]  (.A(\un24_next_sum_m[13] ), .B(
        next_sum_0_sqmuxa_1), .C(\un3_next_sum_m[13] ), .Y(
        \un1_next_sum_iv_2[13] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I210_Y (.A(N695), .B(N688), .C(
        N687), .Y(N769));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I15_G0N (.A(\un1_next_sum[15] )
        , .B(sum_15), .Y(N516));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I425_Y_0 (.A(sum_7), .B(
        \un1_next_sum[7] ), .Y(ADD_40x40_fast_I425_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I139_Y (.A(N611), .B(N615), .Y(
        N692));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I384_un1_Y (.A(N882), .B(N666), 
        .C(N850), .Y(I384_un1_Y));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I277_Y (.A(N706), .B(N698), .C(
        N764), .Y(N848));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I159_Y (.A(N635), .B(N631), .Y(
        N712));
    DFN1E1C0 \i_adj[13]  (.D(\inf_abs2_5[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[13]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I104_Y (.A(N486), .B(N490), .C(
        N489), .Y(N654));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I115_un1_Y (.A(N393), .B(N266), 
        .Y(I115_un1_Y));
    NOR3 inf_abs2_a_0_I_29 (.A(integral[13]), .B(integral[12]), .C(
        integral[14]), .Y(\DWACT_FINC_E[5] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I130_Y_0 (.A(N386), .B(N379), .C(
        N378), .Y(ADD_22x22_fast_I130_Y_0));
    DFN1E1C0 \preg[12]  (.D(\p_adj[6]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[12]_net_1 ));
    MX2 \i_adj_RNO[2]  (.A(integral[8]), .B(\inf_abs2_a_0[2] ), .S(
        integral_0_0), .Y(\inf_abs2_5[2] ));
    DFN1E1C0 \i_adj[5]  (.D(\inf_abs2_5[5] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[5]_net_1 ));
    DFN1E1C0 \ireg[20]  (.D(\next_ireg_3[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[20]_net_1 ));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I379_Y_0 (.A(\sumreg[36]_net_1 )
        , .B(\sumreg[37]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(
        ADD_40x40_fast_I379_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I321_un1_Y (.A(N816), .B(
        \un1_next_sum[0] ), .Y(I321_un1_Y));
    OR3 un1_sumreg_0_0_ADD_m8_i_o4_1 (.A(sum_2_d0), .B(sum_1_d0), .C(
        sum_0_d0), .Y(ADD_m8_i_o4_1));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I378_Y_0 (.A(\sumreg[38]_net_1 )
        , .B(\sumreg[37]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(
        ADD_40x40_fast_I378_Y_0));
    OR2 next_ireg_3_0_ADD_22x22_fast_I2_P0N (.A(\i_adj[2]_net_1 ), .B(
        \i_adj[4]_net_1 ), .Y(N273));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I134_Y (.A(N606), .B(N610), .Y(
        N687));
    DFN1E1C0 \i_adj[0]  (.D(\inf_abs2_5[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[0]_net_1 ));
    DFN1E1C0 \p_adj[6]  (.D(\inf_abs1_5[6] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[6]_net_1 ));
    MX2 \p_adj_RNO[4]  (.A(sr_new[4]), .B(\inf_abs1_a_2[4] ), .S(
        sr_new_0_0), .Y(\inf_abs1_5[4] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I154_Y (.A(N630), .B(N627), .C(
        N626), .Y(N707));
    AO1 \ireg_RNI7U191[16]  (.A(\ireg[16]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[16] ), .Y(
        \un1_next_sum_iv_1[16] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I211_Y (.A(N688), .B(N696), .Y(
        N770));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I12_G0N (.A(\un1_next_sum[12] )
        , .B(sum_12), .Y(N507_0));
    XA1B \sumreg_RNO[24]  (.A(N1058), .B(ADD_40x40_fast_I442_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[24] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I59_Y (.A(N328), .B(N332), .Y(
        N367));
    MX2 \i_adj_RNO[0]  (.A(integral[6]), .B(integral[6]), .S(
        integral_0_0), .Y(\inf_abs2_5[0] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I57_Y (.A(N326), .B(N330), .Y(
        N365));
    AND3 inf_abs2_a_0_I_42 (.A(\DWACT_FINC_E_0[6] ), .B(
        \DWACT_FINC_E_0[7] ), .C(\DWACT_FINC_E[9] ), .Y(N_12_0));
    NOR2B \preg_RNITIAK[16]  (.A(\preg[16]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[16] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I218_Y (.A(N703), .B(N696), .C(
        N695), .Y(N777));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I168_Y_0 (.A(\i_adj[10]_net_1 ), 
        .B(\i_adj[8]_net_1 ), .Y(ADD_22x22_fast_I168_Y_0));
    XNOR2 inf_abs2_a_0_I_23 (.A(integral[14]), .B(N_19), .Y(
        \inf_abs2_a_0[8] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I66_Y (.A(N339), .B(N336), .C(
        N335), .Y(N374));
    AO1 next_ireg_3_0_ADD_22x22_fast_I44_Y (.A(N281), .B(N285), .C(
        N284), .Y(N349));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I439_Y_0 (.A(sum_21), .B(
        \un1_next_sum[21] ), .Y(ADD_40x40_fast_I439_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I450_Y_0 (.A(
        \sumreg[32]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I450_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I234_Y (.A(N719), .B(N712), .C(
        N711), .Y(N793));
    NOR3B \un1_next_sum_iv_0_RNO[21]  (.A(integral_0_0), .B(
        \state_0[3]_net_1 ), .C(\ireg[21]_net_1 ), .Y(
        \un3_next_sum_m[21] ));
    NOR3B \ireg_RNI45KQ[12]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[12]_net_1 ), .Y(\un3_next_sum_m[12] ));
    NOR3 inf_abs1_a_2_I_33 (.A(sr_new[10]), .B(sr_new[9]), .C(
        sr_new[11]), .Y(\DWACT_FINC_E[7] ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I384_Y (.A(N850), .B(N881), .C(
        ADD_40x40_fast_I384_Y_2), .Y(N1033));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I254_Y (.A(I254_un1_Y), .B(N731), 
        .Y(N813));
    MX2 \i_adj_RNO[7]  (.A(integral[13]), .B(\inf_abs2_a_0[7] ), .S(
        integral_0_0), .Y(\inf_abs2_5[7] ));
    DFN1E1C0 \i_adj[21]  (.D(\inf_abs2_5[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[21]_net_1 ));
    XA1B \sumreg_RNO[9]  (.A(N1103), .B(ADD_40x40_fast_I427_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[9] ));
    OR2 \un1_next_sum_iv[19]  (.A(N_228_1), .B(
        \un1_next_sum_iv_0[19]_net_1 ), .Y(\un1_next_sum[19] ));
    AO1B un1_sumreg_0_0_ADD_40x40_fast_I59_Y (.A(\sumreg[29]_net_1 ), 
        .B(\sumreg[28]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N609)
        );
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I162_Y (.A(N638), .B(N635), .C(
        N634), .Y(N715));
    DFN1E1C0 \ireg[14]  (.D(\next_ireg_3[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[14]_net_1 ));
    DFN1E1C0 \p_adj[11]  (.D(\inf_abs1_5[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\p_adj[11]_net_1 ));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I82_Y (.A(N519), .B(sum_17), .C(
        \un1_next_sum[17] ), .Y(N632));
    NOR2A \state_RNITH09_0[5]  (.A(\state[5]_net_1 ), .B(sr_new[12]), 
        .Y(next_sum_1_sqmuxa_2));
    DFN1E1C0 \i_adj[16]  (.D(\inf_abs2_5[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[16]_net_1 ));
    NOR2B \preg_RNIUJAK[17]  (.A(\preg[17]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .Y(\preg_m[17] ));
    OR2 next_ireg_3_0_ADD_22x22_fast_I4_P0N (.A(\i_adj[6]_net_1 ), .B(
        \i_adj[4]_net_1 ), .Y(N279));
    NOR2B \state_RNI13UM[4]  (.A(\state[4]_net_1 ), .B(derivative_0), 
        .Y(next_sum_0_sqmuxa_1));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I437_Y_0 (.A(sum_19), .B(
        \un1_next_sum[19] ), .Y(ADD_40x40_fast_I437_Y_0));
    NOR3B \un1_next_sum_iv_0_RNO[19]  (.A(integral_0_0), .B(
        \state_0[3]_net_1 ), .C(\ireg[19]_net_1 ), .Y(
        \un3_next_sum_m[19] ));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I13_P0N (.A(\un1_next_sum[13] ), 
        .B(sum_13), .Y(N511));
    MAJ3 next_ireg_3_0_ADD_22x22_fast_I32_Y (.A(N299), .B(
        \i_adj[12]_net_1 ), .C(\i_adj[14]_net_1 ), .Y(N337));
    MX2 \i_adj_RNO[11]  (.A(integral[17]), .B(\inf_abs2_a_0[11] ), .S(
        integral_1_0), .Y(\inf_abs2_5[11] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I130_un1_Y_0 (.A(N387), .B(N379)
        , .Y(ADD_22x22_fast_I130_un1_Y_0));
    OR2 \preg_RNI69KC2[6]  (.A(\un3_next_sum_m[6] ), .B(
        \un1_next_sum_iv_0[6] ), .Y(\un1_next_sum_iv_2[6] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I15_G0N (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .Y(N311));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I298_Y (.A(I298_un1_Y), .B(N785), 
        .Y(N869));
    DFN1E1C0 \ireg[4]  (.D(\i_adj[0]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_1[2]_net_1 ), .Q(\ireg[4]_net_1 ));
    MX2 \p_adj_RNO[11]  (.A(sr_new[11]), .B(\inf_abs1_a_2[11] ), .S(
        sr_new[12]), .Y(\inf_abs1_5[11] ));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I172_Y (.A(\i_adj[14]_net_1 ), 
        .B(\i_adj[12]_net_1 ), .C(N510), .Y(\next_ireg_3[18] ));
    XA1B \sumreg_RNO[37]  (.A(N1025), .B(ADD_40x40_fast_I455_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[37] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I381_un1_Y (.A(N876), .B(N823), 
        .C(N844), .Y(I381_un1_Y));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I141_Y (.A(N613), .B(N617), .Y(
        N694));
    AO1A \preg_RNIDMDC1[6]  (.A(\preg[6]_net_1 ), .B(
        next_sum_0_sqmuxa_2), .C(next_sum_0_sqmuxa_1), .Y(
        \un1_next_sum_iv_0[6] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I83_Y (.A(N356), .B(N352), .Y(
        N391));
    NOR2B \state_RNIGPKC[0]  (.A(sum_enable), .B(sum_rdy), .Y(
        \state_RNIGPKC[0]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I111_Y (.A(N393), .B(N385), .Y(
        N425));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I175_Y (.A(N651), .B(N647), .Y(
        N728));
    DFN1E1C0 \sumreg[24]  (.D(\next_sum[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(\sumreg[24]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I26_Y (.A(N308), .B(N312), .C(
        N311), .Y(N331));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I175_Y (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[17]_net_1 ), .C(N501), .Y(\next_ireg_3[21] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I431_Y_0 (.A(sum_13), .B(
        \un1_next_sum[13] ), .Y(ADD_40x40_fast_I431_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I300_Y (.A(N803), .B(N788), .C(
        N787), .Y(N871));
    NOR3B \ireg_RNI37QU[10]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[10]_net_1 ), .C(integral_1_0), .Y(\ireg_m[10] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I103_Y (.A(N493), .B(N490), .Y(
        N653));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I259_un1_Y (.A(N738), .B(N745), 
        .Y(I259_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I88_Y (.A(N510_0), .B(N514), .C(
        N513), .Y(N638));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I0_P0N (.A(N_228), .B(sum_0_d0), 
        .Y(N472));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I260_Y (.A(N740), .B(N666), .C(
        N739), .Y(N821));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I8_P0N (.A(\un1_next_sum[8] ), 
        .B(sum_8), .Y(N496));
    OR2 \ireg_RNIJ3293[17]  (.A(\un1_next_sum_iv_2[17] ), .B(
        \un1_next_sum_iv_1[17] ), .Y(\un1_next_sum[17] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I379_un1_Y_0 (.A(N872), .B(
        N840), .Y(ADD_40x40_fast_I379_un1_Y_0));
    MX2 \i_adj_RNO[15]  (.A(integral[21]), .B(\inf_abs2_a_0[15] ), .S(
        integral_1_0), .Y(\inf_abs2_5[15] ));
    DFN1E1C0 \sumreg[14]  (.D(\next_sum[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_14));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I350_Y (.A(I290_un1_Y), .B(N777), 
        .C(I350_un1_Y), .Y(N1049));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I203_Y (.A(N680), .B(N688), .Y(
        N762));
    NOR2B \i_adj_RNO[20]  (.A(\inf_abs2_a_0[20] ), .B(integral[25]), 
        .Y(\inf_abs2_5[20] ));
    XNOR2 inf_abs1_a_2_I_14 (.A(sr_new[5]), .B(N_9_0), .Y(
        \inf_abs1_a_2[5] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I170_Y_0 (.A(\i_adj[12]_net_1 ), 
        .B(\i_adj[10]_net_1 ), .Y(ADD_22x22_fast_I170_Y_0));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I133_Y (.A(N605), .B(N609), .Y(
        N686));
    OR2A un1_sumreg_0_0_ADD_40x40_fast_I38_P0N (.A(
        \un1_next_sum_1_iv[26] ), .B(\sumreg[38]_net_1 ), .Y(N586));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I215_Y (.A(N692), .B(N700), .Y(
        N774));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I279_Y (.A(N692), .B(N684), .C(
        N782), .Y(N850));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I153_Y (.A(N625), .B(N629), .Y(
        N706));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I79_Y (.A(N348), .B(N352), .Y(
        N387));
    XA1B \sumreg_RNO[30]  (.A(N1040), .B(ADD_40x40_fast_I448_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[30] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I77_Y (.A(N350), .B(N346), .Y(
        N385));
    XNOR2 inf_abs2_a_0_I_9 (.A(integral[9]), .B(N_24), .Y(
        \inf_abs2_a_0[3] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I233_Y (.A(N710), .B(N718), .Y(
        N792));
    XA1B \sumreg_RNO[31]  (.A(N1037), .B(ADD_40x40_fast_I449_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[31] ));
    NOR3 inf_abs2_a_0_I_10 (.A(integral[7]), .B(integral[6]), .C(
        integral[8]), .Y(\DWACT_FINC_E_0[0] ));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I440_Y_0 (.A(sum_22), .B(
        \un1_next_sum[22] ), .Y(ADD_40x40_fast_I440_Y_0));
    AO1 \preg_RNINH5Q1[7]  (.A(\preg[7]_net_1 ), .B(
        next_sum_1_sqmuxa_2), .C(\ireg_m[7] ), .Y(
        \un1_next_sum_iv_1[7] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I253_Y (.A(N738), .B(N730), .Y(
        N812));
    AO1 next_ireg_3_0_ADD_22x22_fast_I52_Y (.A(N269), .B(N273), .C(
        N272), .Y(N357));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I108_Y (.A(N480), .B(N484), .C(
        N483), .Y(N658));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I261_Y (.A(N472), .B(
        \un1_next_sum[0] ), .C(N741), .Y(N823));
    NOR3 \state_RNIAF301[6]  (.A(sum_rdy), .B(\state[6]_net_1 ), .C(
        \state_0[1]_net_1 ), .Y(N_416_0));
    XOR3 next_ireg_3_0_ADD_22x22_fast_I173_Y (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[13]_net_1 ), .C(N507), .Y(\next_ireg_3[19] ));
    NOR2 inf_abs1_a_2_I_15 (.A(sr_new[3]), .B(sr_new[4]), .Y(
        \DWACT_FINC_E_0[1] ));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I83_Y (.A(sum_17), .B(
        \un1_next_sum[17] ), .C(N520), .Y(N633));
    XA1B \sumreg_RNO[25]  (.A(N1055), .B(ADD_40x40_fast_I443_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[25] ));
    DFN1E1C0 \i_adj[11]  (.D(\inf_abs2_5[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state[1]_net_1 ), .Q(\i_adj[11]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I307_Y (.A(N810), .B(N794), .Y(
        N878));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I138_Y (.A(N614), .B(N611), .C(
        N610), .Y(N691));
    DFN1E1C0 \ireg[11]  (.D(\next_ireg_3[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[11]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I311_Y (.A(N814), .B(N798), .Y(
        N882));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I420_Y_0 (.A(sum_2_d0), .B(
        \un1_next_sum[0] ), .Y(ADD_40x40_fast_I420_Y_0));
    DFN1C0 \state[3]  (.D(\state[6]_net_1 ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[3]_net_1 ));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I158_Y (.A(N634), .B(N631), .C(
        N630), .Y(N711));
    XA1 \ireg_RNI35LQ[20]  (.A(integral_0_0), .B(\ireg[20]_net_1 ), .C(
        \state_0[3]_net_1 ), .Y(\un1_next_sum_iv_0[20] ));
    MX2 \i_adj_RNO[17]  (.A(integral[23]), .B(\inf_abs2_a_0[17] ), .S(
        integral[25]), .Y(\inf_abs2_5[17] ));
    DFN1E1C0 \i_adj[1]  (.D(\inf_abs2_5[1] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\i_adj[1]_net_1 ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I80_Y (.A(N353), .B(N350), .C(
        N349), .Y(N388));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I86_Y (.A(N513), .B(N517), .C(
        N516), .Y(N636));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I236_Y (.A(N721), .B(N714), .C(
        N713), .Y(N795));
    DFN1E1C0 \sumreg[3]  (.D(\next_sum[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_416_0), .Q(sum_3));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I358_un1_Y (.A(N878), .B(N743), 
        .Y(I358_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I220_Y (.A(N705), .B(N698), .C(
        N697), .Y(N779));
    OR2 un1_sumreg_0_0_ADD_40x40_fast_I256_Y (.A(I256_un1_Y), .B(N733), 
        .Y(N815));
    DFN1E1C0 \sumreg_1[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(sum_1_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I382_Y_1 (.A(N762), .B(N777), .C(
        ADD_40x40_fast_I382_Y_0), .Y(ADD_40x40_fast_I382_Y_1));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I4_G0N (.A(\i_adj[6]_net_1 ), 
        .B(\i_adj[4]_net_1 ), .Y(N278));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I357_Y (.A(N876), .B(N823), .C(
        N875), .Y(N1070));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I85_Y (.A(N358), .B(N354), .Y(
        N393));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I142_Y (.A(N618), .B(N615), .C(
        N614), .Y(N695));
    DFN1C0 \state_0[1]  (.D(\state_RNIGPKC[0]_net_1 ), .CLK(clk_c), 
        .CLR(n_rst_c), .Q(\state_0[1]_net_1 ));
    NOR3 inf_abs2_a_0_I_50 (.A(integral[22]), .B(integral[21]), .C(
        integral[23]), .Y(\DWACT_FINC_E[12] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I347_un1_Y_0 (.A(N788), .B(
        N772), .Y(ADD_40x40_fast_I347_un1_Y_0));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I3_G0N (.A(\i_adj[5]_net_1 ), 
        .B(\i_adj[3]_net_1 ), .Y(N275));
    XNOR2 inf_abs1_a_2_I_9 (.A(sr_new[3]), .B(N_11_0), .Y(
        \inf_abs1_a_2[3] ));
    XOR2 next_ireg_3_0_ADD_22x22_fast_I171_Y_0 (.A(\i_adj[11]_net_1 ), 
        .B(\i_adj[13]_net_1 ), .Y(ADD_22x22_fast_I171_Y_0));
    NOR3B inf_abs1_a_2_I_16 (.A(\DWACT_FINC_E_0[1] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[5]), .Y(N_8_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I46_Y (.A(N278), .B(N282), .C(
        N281), .Y(N351));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I13_G0N (.A(\i_adj[15]_net_1 ), 
        .B(\i_adj[13]_net_1 ), .Y(N305));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I361_un1_Y (.A(N884), .B(
        \un1_next_sum[0] ), .Y(I361_un1_Y));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I350_un1_Y (.A(N778), .B(N794), 
        .C(N1097), .Y(I350_un1_Y));
    NOR3B \preg_RNIQFAK[13]  (.A(sr_new[12]), .B(\state[5]_net_1 ), .C(
        \preg[13]_net_1 ), .Y(\un24_next_sum_m[13] ));
    VCC VCC_i (.Y(VCC));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I14_G0N (.A(\un1_next_sum[14] )
        , .B(sum_14), .Y(N513));
    MAJ3 un1_sumreg_0_0_ADD_40x40_fast_I116_Y (.A(sum_0_d0), .B(N_228), 
        .C(\un1_next_sum[0] ), .Y(N666));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I50_Y (.A(\sumreg[33]_net_1 ), 
        .B(\sumreg[32]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N600)
        );
    AND3 inf_abs1_a_2_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(
        \DWACT_FINC_E[4] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I6_G0N (.A(\un1_next_sum[6] ), 
        .B(sum_6), .Y(N489));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I385_Y_1 (.A(N768), .B(N783), .C(
        ADD_40x40_fast_I385_Y_0), .Y(ADD_40x40_fast_I385_Y_1));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I309_Y (.A(N812), .B(N796), .Y(
        N880));
    AO1 next_ireg_3_0_ADD_22x22_fast_I130_Y (.A(
        ADD_22x22_fast_I130_un1_Y_0), .B(N394), .C(
        ADD_22x22_fast_I130_Y_0), .Y(N510));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I383_un1_Y (.A(N880), .B(N745), 
        .C(N848), .Y(I383_un1_Y));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I185_Y (.A(N487), .B(N484), .C(
        N661), .Y(N738));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I448_Y_0 (.A(
        \sumreg[30]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I448_Y_0));
    AO1 next_ireg_3_0_ADD_22x22_fast_I129_Y_0 (.A(N384), .B(N377), .C(
        N376), .Y(ADD_22x22_fast_I129_Y_0));
    XA1 \ireg_RNI7QL41[4]  (.A(integral_1_0), .B(\ireg[4]_net_1 ), .C(
        \state[3]_net_1 ), .Y(\un1_next_sum_iv_0[4] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I246_un1_Y (.A(N731), .B(N724), 
        .Y(I246_un1_Y));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I228_Y (.A(N713), .B(N706), .C(
        N705), .Y(N787));
    OR3 \state_RNIFG0J1[4]  (.A(next_sum_1_sqmuxa_2), .B(
        next_sum_1_sqmuxa_1), .C(next_sum_1_sqmuxa), .Y(
        \un1_next_sum_1_iv_0[26] ));
    NOR3B \ireg_RNI23KQ[10]  (.A(integral_0_0), .B(\state_0[3]_net_1 ), 
        .C(\ireg[10]_net_1 ), .Y(\un3_next_sum_m[10] ));
    NOR3 inf_abs1_a_2_I_8 (.A(sr_new[0]), .B(sr_new[2]), .C(sr_new[1]), 
        .Y(N_11_0));
    XA1B \sumreg_RNO[26]  (.A(N1052), .B(ADD_40x40_fast_I444_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[26] ));
    OR2 \ireg_RNI5FK42[4]  (.A(\un1_next_sum_iv_0[4] ), .B(N_228_1), 
        .Y(\un1_next_sum[4] ));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I454_Y_0 (.A(
        \sumreg[36]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I454_Y_0));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I110_Y (.A(sum_2_d0), .B(
        \un1_next_sum[0] ), .C(N480), .Y(N660));
    XA1B \sumreg_RNO[17]  (.A(N1079), .B(ADD_40x40_fast_I435_Y_0), .C(
        \state_2[2]_net_1 ), .Y(\next_sum[17] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I286_un1_Y (.A(N789), .B(N774), 
        .Y(I286_un1_Y));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I359_Y (.A(N795), .B(I308_un1_Y), 
        .C(I359_un1_Y), .Y(N1076));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I137_Y (.A(N613), .B(N609), .Y(
        N690));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I129_un1_Y_0 (.A(N377), .B(N385)
        , .Y(ADD_22x22_fast_I129_un1_Y_0));
    XNOR2 un1_sumreg_0_0_ADD_40x40_fast_I453_Y_0 (.A(
        \sumreg[35]_net_1 ), .B(\un1_next_sum_1_iv[26] ), .Y(
        ADD_40x40_fast_I453_Y_0));
    OA1B un1_sumreg_0_0_ADD_40x40_fast_I48_Y (.A(\sumreg[34]_net_1 ), 
        .B(\sumreg[33]_net_1 ), .C(\un1_next_sum_1_iv_0[26] ), .Y(N598)
        );
    NOR2A inf_abs1_a_2_I_25 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .Y(
        N_5));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I157_Y (.A(N629), .B(N633), .Y(
        N710));
    XOR2 un1_sumreg_0_0_ADD_40x40_fast_I428_Y_0 (.A(sum_10), .B(
        \un1_next_sum[10] ), .Y(ADD_40x40_fast_I428_Y_0));
    DFN1E1C0 \preg[11]  (.D(\p_adj[5]_net_1 ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\preg[11]_net_1 ));
    XA1B \sumreg_RNO[23]  (.A(N1061), .B(ADD_40x40_fast_I441_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[23] ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I131_un1_Y (.A(N421), .B(N396), 
        .Y(I131_un1_Y));
    DFN1E1C0 \sumreg[22]  (.D(\next_sum[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(sum_22));
    OR2 next_ireg_3_0_ADD_22x22_fast_I115_Y (.A(I115_un1_Y), .B(N392), 
        .Y(N531));
    OR3 un1_sumreg_0_0_ADD_40x40_fast_I5_P0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[5] ), .C(sum_5), .Y(N487));
    NOR3B \ireg_RNI48QU[11]  (.A(\state_0[3]_net_1 ), .B(
        \ireg[11]_net_1 ), .C(integral_1_0), .Y(\ireg_m[11] ));
    NOR3C un1_sumreg_0_0_ADD_40x40_fast_I66_un1_Y (.A(
        \sumreg[24]_net_1 ), .B(\un1_next_sum[24] ), .C(N547), .Y(
        I66_un1_Y));
    OA1 un1_sumreg_0_0_ADD_40x40_fast_I20_G0N (.A(N_228_1), .B(
        \un1_next_sum_iv_0[20] ), .C(sum_20), .Y(N531_0));
    DFN1E1C0 \ireg[13]  (.D(\next_ireg_3[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[13]_net_1 ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I296_un1_Y (.A(N799), .B(N784), 
        .Y(I296_un1_Y));
    XA1B \sumreg_RNO[29]  (.A(N1043), .B(ADD_40x40_fast_I447_Y_0), .C(
        \state[2]_net_1 ), .Y(\next_sum[29] ));
    NOR2A \state_RNI13UM_0[4]  (.A(\state[4]_net_1 ), .B(derivative_0), 
        .Y(next_sum_1_sqmuxa_1));
    DFN1E1C0 \p_adj[8]  (.D(\inf_abs1_5[8] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[1]_net_1 ), .Q(\p_adj[8]_net_1 ));
    NOR2B next_ireg_3_0_ADD_22x22_fast_I61_Y (.A(N334), .B(N330), .Y(
        N369));
    AX1D next_ireg_3_0_ADD_22x22_fast_I177_Y (.A(I124_un1_Y), .B(
        ADD_22x22_fast_I144_Y_2), .C(ADD_22x22_fast_I177_Y_0), .Y(
        \next_ireg_3[23] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I84_Y (.A(N357), .B(N354), .C(
        N353), .Y(N392));
    AO1 un1_sumreg_0_0_ADD_40x40_fast_I240_Y (.A(N725), .B(N718), .C(
        N717), .Y(N799));
    XNOR2 inf_abs1_a_2_I_7 (.A(sr_new[2]), .B(N_12), .Y(
        \inf_abs1_a_2[2] ));
    XNOR2 inf_abs2_a_0_I_17 (.A(integral[12]), .B(N_21), .Y(
        \inf_abs2_a_0[6] ));
    DFN1E1C0 \sumreg[12]  (.D(\next_sum[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416_0), .Q(sum_12));
    DFN1E1C0 \ireg[15]  (.D(\next_ireg_3[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(\state_0[2]_net_1 ), .Q(\ireg[15]_net_1 ));
    XA1B \sumreg_RNO[1]  (.A(N666), .B(ADD_40x40_fast_I419_Y_0), .C(
        \state_1[2]_net_1 ), .Y(\next_sum[1] ));
    AO1 next_ireg_3_0_ADD_22x22_fast_I72_Y (.A(N345), .B(N342), .C(
        N341), .Y(N380));
    AX1D next_ireg_3_0_ADD_22x22_fast_I179_Y (.A(I120_un1_Y), .B(
        ADD_22x22_fast_I142_Y_3), .C(ADD_22x22_fast_I179_Y_0), .Y(
        \next_ireg_3[25] ));
    NOR2B un1_sumreg_0_0_ADD_40x40_fast_I97_Y (.A(N502), .B(N499), .Y(
        N647));
    OR2 next_ireg_3_0_ADD_22x22_fast_I8_P0N (.A(\i_adj[8]_net_1 ), .B(
        \i_adj[10]_net_1 ), .Y(N291));
    DFN1E1C0 \sumreg_2[39]  (.D(\next_sum[39] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_416), .Q(sum_2_0));
    OR2 \preg_RNIVSP64[7]  (.A(\un1_next_sum_iv_2[7] ), .B(
        \un1_next_sum_iv_1[7] ), .Y(\un1_next_sum[7] ));
    AO1 \ireg_RNIB2291[18]  (.A(\ireg[18]_net_1 ), .B(
        next_sum_1_sqmuxa), .C(\preg_m[18] ), .Y(
        \un1_next_sum_iv_1[18] ));
    NOR3 inf_abs1_a_2_I_18 (.A(sr_new[4]), .B(sr_new[3]), .C(sr_new[5])
        , .Y(\DWACT_FINC_E_0[2] ));
    XNOR2 inf_abs1_a_2_I_26 (.A(sr_new[9]), .B(N_5), .Y(
        \inf_abs1_a_2[9] ));
    
endmodule


module sig_gen_7(
       vd_done,
       n_rst_c,
       clk_c,
       sig_old_i_0,
       sig_prev
    );
input  vd_done;
input  n_rst_c;
input  clk_c;
output sig_old_i_0;
output sig_prev;

    wire sig_prev_i, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(clk_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev_inst_1 (.D(vd_done), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(sig_prev));
    INV sig_old_RNO (.A(sig_prev), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module spi_stp_12s_1_4(
       cur_vd,
       N_29,
       din_15_c,
       n_rst_c,
       sck_5_c
    );
output [11:0] cur_vd;
input  N_29;
input  din_15_c;
input  n_rst_c;
input  sck_5_c;

    wire GND, VCC;
    
    DFN1E0C0 \sr[7]  (.D(cur_vd[6]), .CLK(sck_5_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[7]));
    DFN1E0C0 \sr[5]  (.D(cur_vd[4]), .CLK(sck_5_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[5]));
    DFN1E0C0 \sr[10]  (.D(cur_vd[9]), .CLK(sck_5_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[10]));
    DFN1E0C0 \sr[8]  (.D(cur_vd[7]), .CLK(sck_5_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[8]));
    DFN1E0C0 \sr[3]  (.D(cur_vd[2]), .CLK(sck_5_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[3]));
    DFN1E0C0 \sr[1]  (.D(cur_vd[0]), .CLK(sck_5_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[1]));
    DFN1E0C0 \sr[2]  (.D(cur_vd[1]), .CLK(sck_5_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[2]));
    DFN1E0C0 \sr[9]  (.D(cur_vd[8]), .CLK(sck_5_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[9]));
    VCC VCC_i (.Y(VCC));
    DFN1E0C0 \sr[11]  (.D(cur_vd[10]), .CLK(sck_5_c), .CLR(n_rst_c), 
        .E(N_29), .Q(cur_vd[11]));
    DFN1E0C0 \sr[0]  (.D(din_15_c), .CLK(sck_5_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[0]));
    GND GND_i (.Y(GND));
    DFN1E0C0 \sr[6]  (.D(cur_vd[5]), .CLK(sck_5_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[6]));
    DFN1E0C0 \sr[4]  (.D(cur_vd[3]), .CLK(sck_5_c), .CLR(n_rst_c), .E(
        N_29), .Q(cur_vd[4]));
    
endmodule


module sig_gen_0_1(
       cs_i_1,
       n_rst_c,
       sck_5_c,
       vd_done
    );
input  cs_i_1;
input  n_rst_c;
input  sck_5_c;
output vd_done;

    wire sig_prev_i, sig_prev_net_1, sig_old_i_0, GND, VCC;
    
    VCC VCC_i (.Y(VCC));
    NOR2B sig_old_RNIAHVF (.A(sig_prev_net_1), .B(sig_old_i_0), .Y(
        vd_done));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(sck_5_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev (.D(cs_i_1), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        sig_prev_net_1));
    INV sig_old_RNO (.A(sig_prev_net_1), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module spi_ctl_12s_2(
       n_rst_c,
       sck_5_c,
       N_29,
       cs_i_1,
       cs_i_1_i
    );
input  n_rst_c;
input  sck_5_c;
output N_29;
output cs_i_1;
output cs_i_1_i;

    wire cnt_m1_0_a2_0, \cnt[14]_net_1 , \cnt[13]_net_1 , 
        cnt_m6_0_a2_6, cnt_m6_0_a2_0, \cnt[3]_net_1 , cnt_m5_0_a2_2, 
        cnt_m6_0_a2_2, \cnt[7]_net_1 , \cnt[8]_net_1 , \cnt[11]_net_1 , 
        \cnt[10]_net_1 , cnt_m7_0_a2_4, \cnt[5]_net_1 , cnt_m7_0_a2_3, 
        \cnt[6]_net_1 , cnt_m7_0_a2_1, \cnt[9]_net_1 , 
        state_tr0_0_a3_12, state_tr0_0_a3_6, state_tr0_0_a3_9, N_103, 
        \cnt[4]_net_1 , state_tr0_0_a3_8, state_tr0_0_a3_4, 
        state_tr0_0_a3_7, state_tr0_0_a3_2, \cnt[0]_net_1 , 
        \cnt[1]_net_1 , state_tr0_0_a3_1, \cnt[15]_net_1 , 
        \cnt[12]_net_1 , vd_stp_en_i_a3_9, vd_stp_en_i_a3_4, 
        vd_stp_en_i_a3_3, N_73, vd_stp_en_i_a3_8, vd_stp_en_i_a3_2, 
        vd_stp_en_i_a3_5, cnt_m6_0_a2_5_6, cnt_m6_0_a2_5_0, 
        cnt_m6_0_a2_5, \cnt[2]_net_1 , cnt_m5_0_a2_3, cnt_m2_0_a2_0, 
        cnt_m5_0_a2_1, cnt_m2_0_a2_2, cnt_m2_0_a2_1, N_74, 
        cnt_N_13_mux, N_33, N_31, cnt_N_7_mux_0_0, cnt_N_3_mux_0, 
        cnt_N_11_mux_2, cnt_N_15_mux, cnt_N_13_mux_0, N_30, 
        \state_RNO_8[0] , N_26, N_24, N_22, N_20, N_97, N_18, N_14, 
        N_12, N_36, \cnt_RNO[6]_net_1 , cnt_n10, d_N_3_mux, 
        \cnt_RNO_1_3[10] , cnt_n0, cnt_n15, cnt_n14, cnt_n13, N_72, 
        cnt_n12, cnt_n11, cnt_n9, N_38, GND, VCC;
    
    NOR2B \cnt_RNO_2[6]  (.A(\cnt[4]_net_1 ), .B(\cnt[3]_net_1 ), .Y(
        cnt_m2_0_a2_2));
    XA1A \cnt_RNO[8]  (.A(\cnt[8]_net_1 ), .B(N_36), .C(cs_i_1), .Y(
        N_12));
    NOR2 \cnt_RNIOVKI[9]  (.A(\cnt[9]_net_1 ), .B(\cnt[7]_net_1 ), .Y(
        vd_stp_en_i_a3_4));
    NOR2 \cnt_RNIDKKI[2]  (.A(\cnt[3]_net_1 ), .B(\cnt[2]_net_1 ), .Y(
        N_103));
    NOR3C \cnt_RNO_3[10]  (.A(\cnt[3]_net_1 ), .B(\cnt[5]_net_1 ), .C(
        cs_i_1), .Y(cnt_m7_0_a2_4));
    NOR3B \cnt_RNI00B43[3]  (.A(cnt_m6_0_a2_6), .B(cnt_m6_0_a2_5), .C(
        N_31), .Y(cnt_N_13_mux));
    NOR3A \state_RNO_0[0]  (.A(state_tr0_0_a3_4), .B(\cnt[6]_net_1 ), 
        .C(\cnt[7]_net_1 ), .Y(state_tr0_0_a3_8));
    XA1A \cnt_RNO[2]  (.A(N_30), .B(\cnt[2]_net_1 ), .C(cs_i_1), .Y(
        N_24));
    AO1B \state_RNI91L93[0]  (.A(vd_stp_en_i_a3_9), .B(
        vd_stp_en_i_a3_8), .C(cs_i_1), .Y(N_29));
    DFN1C0 \cnt[2]  (.D(N_24), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[2]_net_1 ));
    DFN1C0 \cnt[8]  (.D(N_12), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[8]_net_1 ));
    DFN1C0 \cnt[1]  (.D(N_26), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[1]_net_1 ));
    OA1C \cnt_RNO_0[4]  (.A(\cnt[3]_net_1 ), .B(N_31), .C(
        \cnt[4]_net_1 ), .Y(N_97));
    NOR3C \cnt_RNIJ8231[3]  (.A(cnt_m6_0_a2_0), .B(\cnt[3]_net_1 ), .C(
        cnt_m5_0_a2_2), .Y(cnt_m6_0_a2_6));
    DFN1C0 \cnt[11]  (.D(cnt_n11), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[11]_net_1 ));
    NOR3C \cnt_RNO_0[6]  (.A(cnt_m2_0_a2_1), .B(cnt_m2_0_a2_0), .C(
        cnt_m2_0_a2_2), .Y(cnt_N_7_mux_0_0));
    NOR2B \cnt_RNO_1[15]  (.A(\cnt[14]_net_1 ), .B(\cnt[13]_net_1 ), 
        .Y(cnt_m1_0_a2_0));
    XA1A \cnt_RNO[3]  (.A(N_31), .B(\cnt[3]_net_1 ), .C(cs_i_1), .Y(
        N_22));
    OR2B \cnt_RNO_0[13]  (.A(cnt_N_13_mux), .B(\cnt[12]_net_1 ), .Y(
        N_72));
    NOR3B \state_RNO_6[0]  (.A(\cnt[5]_net_1 ), .B(N_103), .C(
        \cnt[4]_net_1 ), .Y(state_tr0_0_a3_9));
    VCC VCC_i (.Y(VCC));
    NOR2B \cnt_RNI9GKI_0[1]  (.A(\cnt[1]_net_1 ), .B(\cnt[0]_net_1 ), 
        .Y(cnt_m2_0_a2_0));
    XA1 \cnt_RNO[1]  (.A(\cnt[0]_net_1 ), .B(\cnt[1]_net_1 ), .C(
        cs_i_1), .Y(N_26));
    OR2A \cnt_RNI50VR[4]  (.A(\cnt[4]_net_1 ), .B(N_103), .Y(N_73));
    DFN1C0 \cnt[6]  (.D(\cnt_RNO[6]_net_1 ), .CLK(sck_5_c), .CLR(
        n_rst_c), .Q(\cnt[6]_net_1 ));
    NOR3C \cnt_RNO_0[15]  (.A(cnt_m1_0_a2_0), .B(\cnt[12]_net_1 ), .C(
        cnt_N_13_mux), .Y(cnt_N_3_mux_0));
    OR2B \cnt_RNISPIA2[7]  (.A(cnt_N_11_mux_2), .B(\cnt[7]_net_1 ), .Y(
        N_36));
    NOR3A \state_RNO_1[0]  (.A(state_tr0_0_a3_2), .B(\cnt[0]_net_1 ), 
        .C(\cnt[1]_net_1 ), .Y(state_tr0_0_a3_7));
    DFN1C0 \cnt[4]  (.D(N_20), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[4]_net_1 ));
    DFN1C0 \cnt[9]  (.D(cnt_n9), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[9]_net_1 ));
    NOR2A \cnt_RNO[0]  (.A(cs_i_1), .B(\cnt[0]_net_1 ), .Y(cnt_n0));
    OR3C \cnt_RNO_0[14]  (.A(\cnt[12]_net_1 ), .B(\cnt[13]_net_1 ), .C(
        cnt_N_13_mux), .Y(N_74));
    DFN1C0 \cnt[0]  (.D(cnt_n0), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[0]_net_1 ));
    NOR3B \cnt_RNO[4]  (.A(N_33), .B(cs_i_1), .C(N_97), .Y(N_20));
    NOR3 \cnt_RNICQDG[15]  (.A(\cnt[14]_net_1 ), .B(\cnt[15]_net_1 ), 
        .C(\cnt[5]_net_1 ), .Y(vd_stp_en_i_a3_5));
    NOR3C \cnt_RNI69KU[10]  (.A(vd_stp_en_i_a3_2), .B(state_tr0_0_a3_1)
        , .C(vd_stp_en_i_a3_5), .Y(vd_stp_en_i_a3_8));
    NOR2 \state_RNO_4[0]  (.A(\cnt[10]_net_1 ), .B(\cnt[8]_net_1 ), .Y(
        state_tr0_0_a3_2));
    NOR2B \cnt_RNIGNKI[2]  (.A(\cnt[2]_net_1 ), .B(\cnt[6]_net_1 ), .Y(
        cnt_m5_0_a2_1));
    OR3B \cnt_RNIEGJE1[4]  (.A(\cnt[3]_net_1 ), .B(\cnt[4]_net_1 ), .C(
        N_31), .Y(N_33));
    DFN1C0 \state[0]  (.D(\state_RNO_8[0] ), .CLK(sck_5_c), .CLR(
        n_rst_c), .Q(cs_i_1));
    XA1 \cnt_RNO[6]  (.A(cnt_N_7_mux_0_0), .B(\cnt[6]_net_1 ), .C(
        cs_i_1), .Y(\cnt_RNO[6]_net_1 ));
    XA1 \cnt_RNO[15]  (.A(\cnt[15]_net_1 ), .B(cnt_N_3_mux_0), .C(
        cs_i_1), .Y(cnt_n15));
    XA1A \cnt_RNO[9]  (.A(\cnt[9]_net_1 ), .B(N_38), .C(cs_i_1), .Y(
        cnt_n9));
    GND GND_i (.Y(GND));
    NOR2B \cnt_RNO_5[10]  (.A(\cnt[8]_net_1 ), .B(\cnt[9]_net_1 ), .Y(
        cnt_m7_0_a2_1));
    NOR3C \cnt_RNIET951[9]  (.A(\cnt[9]_net_1 ), .B(\cnt[6]_net_1 ), 
        .C(cnt_m6_0_a2_2), .Y(cnt_m6_0_a2_5));
    NOR2B \cnt_RNIB537[11]  (.A(\cnt[11]_net_1 ), .B(\cnt[10]_net_1 ), 
        .Y(cnt_m6_0_a2_0));
    DFN1C0 \cnt[13]  (.D(cnt_n13), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[13]_net_1 ));
    NOR3A \state_RNO_5[0]  (.A(state_tr0_0_a3_1), .B(\cnt[14]_net_1 ), 
        .C(\cnt[15]_net_1 ), .Y(state_tr0_0_a3_6));
    OR2B \cnt_RNI9GKI[1]  (.A(\cnt[1]_net_1 ), .B(\cnt[0]_net_1 ), .Y(
        N_30));
    OR2A \cnt_RNO_0[9]  (.A(\cnt[8]_net_1 ), .B(N_36), .Y(N_38));
    DFN1C0 \cnt[7]  (.D(N_14), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[7]_net_1 ));
    NOR3C \state_RNO_2[0]  (.A(state_tr0_0_a3_6), .B(cs_i_1), .C(
        state_tr0_0_a3_9), .Y(state_tr0_0_a3_12));
    DFN1C0 \cnt[10]  (.D(cnt_n10), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[10]_net_1 ));
    NOR3C \cnt_RNO_1[11]  (.A(cnt_m6_0_a2_5_0), .B(\cnt[3]_net_1 ), .C(
        cnt_m5_0_a2_2), .Y(cnt_m6_0_a2_5_6));
    XA1A \cnt_RNO[5]  (.A(\cnt[5]_net_1 ), .B(N_33), .C(cs_i_1), .Y(
        N_18));
    NOR2 \cnt_RNIE837[11]  (.A(\cnt[11]_net_1 ), .B(\cnt[13]_net_1 ), 
        .Y(state_tr0_0_a3_1));
    NOR3C \cnt_RNI1B812[2]  (.A(cnt_m5_0_a2_2), .B(cnt_m5_0_a2_1), .C(
        cnt_m5_0_a2_3), .Y(cnt_N_11_mux_2));
    DFN1C0 \cnt[3]  (.D(N_22), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[3]_net_1 ));
    NOR2B \cnt_RNO_2[11]  (.A(\cnt[10]_net_1 ), .B(\cnt[2]_net_1 ), .Y(
        cnt_m6_0_a2_5_0));
    XA1A \cnt_RNO[14]  (.A(\cnt[14]_net_1 ), .B(N_74), .C(cs_i_1), .Y(
        cnt_n14));
    NOR2B \cnt_RNINUKI[7]  (.A(\cnt[7]_net_1 ), .B(\cnt[8]_net_1 ), .Y(
        cnt_m6_0_a2_2));
    XNOR2 \cnt_RNO_1[10]  (.A(\cnt[10]_net_1 ), .B(\cnt[4]_net_1 ), .Y(
        \cnt_RNO_1_3[10] ));
    NOR2 \cnt_RNIMTKI[6]  (.A(\cnt[8]_net_1 ), .B(\cnt[6]_net_1 ), .Y(
        vd_stp_en_i_a3_3));
    OR2A \cnt_RNIVPUR[2]  (.A(\cnt[2]_net_1 ), .B(N_30), .Y(N_31));
    NOR3C \cnt_RNO_4[10]  (.A(\cnt[7]_net_1 ), .B(\cnt[6]_net_1 ), .C(
        cnt_m7_0_a2_1), .Y(cnt_m7_0_a2_3));
    NOR3B \cnt_RNO_0[11]  (.A(cnt_m6_0_a2_5), .B(cnt_m6_0_a2_5_6), .C(
        N_30), .Y(cnt_N_13_mux_0));
    XA1 \cnt_RNO[11]  (.A(\cnt[11]_net_1 ), .B(cnt_N_13_mux_0), .C(
        cs_i_1), .Y(cnt_n11));
    NOR3C \cnt_RNIJT812[4]  (.A(vd_stp_en_i_a3_4), .B(vd_stp_en_i_a3_3)
        , .C(N_73), .Y(vd_stp_en_i_a3_9));
    NOR3B \cnt_RNO_2[10]  (.A(cnt_m7_0_a2_4), .B(cnt_m7_0_a2_3), .C(
        N_31), .Y(cnt_N_15_mux));
    OR3C \state_RNO[0]  (.A(state_tr0_0_a3_8), .B(state_tr0_0_a3_7), 
        .C(state_tr0_0_a3_12), .Y(\state_RNO_8[0] ));
    MX2B \cnt_RNO[10]  (.A(d_N_3_mux), .B(\cnt_RNO_1_3[10] ), .S(
        cnt_N_15_mux), .Y(cnt_n10));
    DFN1C0 \cnt[15]  (.D(cnt_n15), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[15]_net_1 ));
    INV \state_RNIGQN9[0]  (.A(cs_i_1), .Y(cs_i_1_i));
    NOR2B \cnt_RNO_1[6]  (.A(\cnt[2]_net_1 ), .B(\cnt[5]_net_1 ), .Y(
        cnt_m2_0_a2_1));
    NOR2B \cnt_RNIHOKI[5]  (.A(\cnt[4]_net_1 ), .B(\cnt[5]_net_1 ), .Y(
        cnt_m5_0_a2_2));
    NOR2B \cnt_RNO_0[10]  (.A(\cnt[10]_net_1 ), .B(cs_i_1), .Y(
        d_N_3_mux));
    NOR2 \state_RNO_3[0]  (.A(\cnt[9]_net_1 ), .B(\cnt[12]_net_1 ), .Y(
        state_tr0_0_a3_4));
    NOR2B \cnt_RNI0RUR[3]  (.A(\cnt[3]_net_1 ), .B(cnt_m2_0_a2_0), .Y(
        cnt_m5_0_a2_3));
    DFN1C0 \cnt[5]  (.D(N_18), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[5]_net_1 ));
    XA1A \cnt_RNO[13]  (.A(\cnt[13]_net_1 ), .B(N_72), .C(cs_i_1), .Y(
        cnt_n13));
    NOR2 \cnt_RNIC637[10]  (.A(\cnt[10]_net_1 ), .B(\cnt[12]_net_1 ), 
        .Y(vd_stp_en_i_a3_2));
    XA1 \cnt_RNO[12]  (.A(\cnt[12]_net_1 ), .B(cnt_N_13_mux), .C(
        cs_i_1), .Y(cnt_n12));
    DFN1C0 \cnt[12]  (.D(cnt_n12), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[12]_net_1 ));
    XA1 \cnt_RNO[7]  (.A(\cnt[7]_net_1 ), .B(cnt_N_11_mux_2), .C(
        cs_i_1), .Y(N_14));
    DFN1C0 \cnt[14]  (.D(cnt_n14), .CLK(sck_5_c), .CLR(n_rst_c), .Q(
        \cnt[14]_net_1 ));
    
endmodule


module spi_rx_12s_3_1(
       cur_vd,
       vd_done,
       cs_i_1_i,
       sck_5_c,
       n_rst_c,
       din_15_c
    );
output [11:0] cur_vd;
output vd_done;
output cs_i_1_i;
input  sck_5_c;
input  n_rst_c;
input  din_15_c;

    wire N_29, cs_i_1, GND, VCC;
    
    spi_stp_12s_1_4 VD_STP (.cur_vd({cur_vd[11], cur_vd[10], cur_vd[9], 
        cur_vd[8], cur_vd[7], cur_vd[6], cur_vd[5], cur_vd[4], 
        cur_vd[3], cur_vd[2], cur_vd[1], cur_vd[0]}), .N_29(N_29), 
        .din_15_c(din_15_c), .n_rst_c(n_rst_c), .sck_5_c(sck_5_c));
    sig_gen_0_1 SPI_RDYSIG (.cs_i_1(cs_i_1), .n_rst_c(n_rst_c), 
        .sck_5_c(sck_5_c), .vd_done(vd_done));
    VCC VCC_i (.Y(VCC));
    spi_ctl_12s_2 SPICTL (.n_rst_c(n_rst_c), .sck_5_c(sck_5_c), .N_29(
        N_29), .cs_i_1(cs_i_1), .cs_i_1_i(cs_i_1_i));
    GND GND_i (.Y(GND));
    
endmodule


module integral_calc_13s_0_4_3(
       sr_new,
       sr_old,
       sr_new_0_0,
       integral,
       integral_i,
       integral_0_0,
       integral_1_0,
       calc_int,
       N_46_1,
       n_rst_c,
       clk_c
    );
input  [12:0] sr_new;
input  [12:0] sr_old;
input  sr_new_0_0;
output [25:6] integral;
output [25:24] integral_i;
output integral_0_0;
output integral_1_0;
input  calc_int;
output N_46_1;
input  n_rst_c;
input  clk_c;

    wire \un1_integ[25] , N_46_1_0, \state[0]_net_1 , \state[1]_net_1 , 
        \un1_next_int_0_iv_0[13] , next_int_1_sqmuxa, 
        next_int_0_sqmuxa_1, N_12, N_10, \DWACT_FINC_E[0] , N_5, 
        \DWACT_FINC_E[4] , N_2, \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , 
        N_12_0, N_10_0, \DWACT_FINC_E_0[0] , N_5_0, 
        \DWACT_FINC_E_0[4] , N_2_0, \DWACT_FINC_E_0[7] , 
        \DWACT_FINC_E_0[6] , \un1_integ[8] , N658, 
        ADD_26x26_fast_I238_Y_0, \un1_integ[11] , N649, 
        ADD_26x26_fast_I241_Y_0, N529, I192_un1_Y, N535, I195_un1_Y, 
        \un1_next_int[11] , \un1_next_int[8] , ADD_26x26_fast_I255_Y_0, 
        \un1_next_int_0_iv[13] , ADD_26x26_fast_I253_Y_0, 
        ADD_26x26_fast_I252_Y_0, ADD_26x26_fast_I249_Y_0, 
        ADD_26x26_fast_I204_Y_3, N502, N517, ADD_26x26_fast_I204_Y_2, 
        N398, ADD_26x26_fast_I204_Y_0, N455, ADD_26x26_fast_I205_Y_2, 
        N400, ADD_26x26_fast_I205_Y_0, N457, ADD_26x26_fast_I250_Y_0, 
        ADD_26x26_fast_I251_Y_0, ADD_26x26_fast_I248_Y_0, 
        ADD_26x26_fast_I206_Y_2, ADD_26x26_fast_I206_un1_Y_0, N522, 
        ADD_26x26_fast_I206_Y_1, N402, N459, ADD_26x26_fast_I207_Y_2, 
        ADD_26x26_fast_I207_un1_Y_0, N524, ADD_26x26_fast_I207_Y_1, 
        N404, N461, ADD_26x26_fast_I210_Y_1, I136_un1_Y, I180_un1_Y, 
        ADD_26x26_fast_I244_Y_0, ADD_26x26_fast_I243_Y_0, 
        ADD_26x26_fast_I242_Y_0, \un2_next_int_m[12] , 
        \un1_next_int_iv_0[12] , ADD_26x26_fast_I208_Y_1, 
        ADD_26x26_fast_I208_un1_Y_0, N526, ADD_26x26_fast_I208_Y_0, 
        N463, ADD_26x26_fast_I209_Y_1, ADD_26x26_fast_I209_un1_Y_0, 
        N528, ADD_26x26_fast_I209_Y_0, N465, N458, 
        ADD_26x26_fast_I211_Y_0, N469, N462, 
        ADD_26x26_fast_I205_un1_Y_0, N466, N474, N504, 
        ADD_26x26_fast_I213_un1_Y_0, N482, N490, \un1_next_int[0] , 
        ADD_26x26_fast_I240_Y_0, \un1_next_int[10] , 
        ADD_26x26_fast_I211_Y_1_0, N470, N483, I160_un1_Y, N506, N489, 
        I163_un1_Y, N512, N487, I162_un1_Y, N510, N508, N539, 
        ADD_26x26_fast_I237_Y_0, \un1_next_int[7] , 
        ADD_26x26_fast_I235_Y_0, \un2_next_int_m[5] , 
        \un1_next_int_iv_1[5] , \integ[5]_net_1 , 
        ADD_26x26_fast_I234_Y_0, \integ[4]_net_1 , \un1_next_int[4] , 
        ADD_26x26_fast_I233_Y_0, \un1_next_int_iv_0[3] , 
        \un1_next_int_iv_1[3] , \integ[3]_net_1 , 
        ADD_26x26_fast_I232_Y_0, \integ[2]_net_1 , \un1_next_int[2] , 
        ADD_26x26_fast_I127_Y_0, ADD_26x26_fast_I125_Y_0, 
        ADD_26x26_fast_I231_Y_0, \un1_next_int_iv_0[1] , 
        \un1_next_int_iv_1[1] , \integ[1]_net_1 , 
        \un1_next_int_iv_1[11] , \un1_next_int_iv_0[11] , 
        \inf_abs0_m[11] , \inf_abs1[11]_net_1 , 
        \un1_next_int_iv_1[10] , \un1_next_int_iv_0[10] , 
        \inf_abs0_m[10] , \un18_next_int_m[10] , \inf_abs1_m[10] , 
        \inf_abs1_a_1[12] , \un1_next_int_iv_0[7] , 
        \inf_abs1[7]_net_1 , ADD_26x26_fast_I230_Y_0, \integ[0]_net_1 , 
        N_3, \un1_next_int_iv_1[9] , \inf_abs0_m[9] , 
        \un18_next_int_m[9] , \inf_abs1_m[9] , \un1_next_int_iv_1[8] , 
        \inf_abs0_m[8] , \un18_next_int_m[8] , \un2_next_int_m[8] , 
        \un1_next_int_iv_1[6] , \un1_next_int_iv_0[6] , 
        \un2_next_int_m[6] , \un18_next_int_m[6] , \inf_abs0_m[6] , 
        \un1_next_int_iv_1[4] , \un1_next_int_iv_0[4] , 
        \un2_next_int_m[4] , \un18_next_int_m[4] , \inf_abs0_m[4] , 
        \un1_next_int_iv_1[0] , \un2_next_int_m[0] , 
        \un1_next_int_iv_0[0] , \inf_abs1[0]_net_1 , \inf_abs0_m[5] , 
        \un18_next_int_m[5] , \inf_abs1_m[5] , \un2_next_int_m[3] , 
        \inf_abs1[3]_net_1 , \un18_next_int_m[3] , 
        \un1_next_int_iv_1[2] , \inf_abs0[2]_net_1 , 
        \un1_next_int_iv_0[2] , \inf_abs1[2]_net_1 , 
        next_int_1_sqmuxa_1, \inf_abs1_m[2] , \inf_abs0[1]_net_1 , 
        \inf_abs1[1]_net_1 , ADD_26x26_fast_I211_Y_1, 
        ADD_26x26_fast_I211_un1_Y_0, N531, \un1_integ[2] , N493, 
        \un1_integ[12] , N527, I191_un1_Y, I210_un1_Y, N530, N491, 
        N514, I213_un1_Y, N635, I186_un1_Y, N519, \inf_abs1_m[8] , 
        \un1_next_int[6] , \inf_abs1_m[6] , \inf_abs1_m[4] , 
        \un1_integ[19] , \un1_integ[16] , \un1_integ[0] , 
        \un1_integ[4] , \un1_integ[6] , \un1_integ[14] , N523, 
        I189_un1_Y, \un1_integ[5] , \un1_integ[21] , I176_un1_Y, 
        \un1_integ[15] , N637, \un1_integ[13] , N525, I190_un1_Y, 
        \un1_integ[3] , \un1_integ[20] , I178_un1_Y, \un1_integ[22] , 
        I174_un1_Y, N401, N405, \un1_next_int[9] , \un2_next_int_m[9] , 
        I204_un1_Y, N518, N655, \un1_integ[9] , \un1_integ[1] , N442, 
        \un1_integ[7] , \un1_integ[10] , I193_un1_Y, \un1_integ[17] , 
        N633, \un1_integ[18] , \un1_integ[23] , I172_un1_Y, 
        \un1_integ[24] , N619, \inf_abs0_m[7] , \un2_next_int_m[7] , 
        \un2_next_int_m[10] , \un2_next_int_m[11] , I184_un1_Y, 
        I212_un1_Y, N534, I170_un1_Y, I205_un1_Y, N403, N399, N460, 
        N456, N478, N486, I56_un1_Y, N345, N424, N344, N425, N342, 
        I58_un1_Y, N426, N427, I102_un1_Y, N348, N351, N473, N420, 
        N476, N423, I106_un1_Y, N428, N477, I108_un1_Y, N430, N479, 
        N480, N431, N434, N484, N435, N419, N415, N475, N422, 
        I54_un1_Y, N347, N440, N317, N321, N320, N441, N318, N350, 
        N438, N324, N323, N439, I74_un1_Y, N472, N488, I120_un1_Y, 
        N464, I148_un1_Y, N471, I156_un1_Y, N467, I144_un1_Y, 
        I188_un1_Y, I194_un1_Y, \inf_abs0[7]_net_1 , 
        \inf_abs0[10]_net_1 , \inf_abs0[11]_net_1 , \inf_abs0_a_0[7] , 
        \inf_abs0_a_0[10] , \inf_abs0_a_0[11] , \inf_abs1_a_1[7] , 
        \inf_abs1_a_1[11] , \inf_abs0_a_0[1] , \inf_abs1_a_1[1] , 
        \inf_abs1_a_1[10] , \inf_abs1_a_1[9] , \inf_abs0_a_0[9] , 
        \inf_abs1_a_1[5] , \inf_abs0_a_0[5] , N417, N416, N413, N406, 
        N407, N408, N409, N412, I146_un1_Y, N410, N411, N414, N485, 
        N418, I96_un1_Y, I50_un1_Y, N353, N354, \inf_abs1[8]_net_1 , 
        \inf_abs1_a_1[8] , \inf_abs1[6]_net_1 , \inf_abs1_a_1[6] , 
        \inf_abs1[4]_net_1 , \inf_abs1_a_1[4] , \inf_abs1_a_1[3] , 
        \inf_abs0_a_0[8] , \inf_abs0_a_0[6] , \inf_abs0_a_0[4] , 
        \inf_abs0_a_0[3] , I142_un1_Y, N336, N481, I150_un1_Y, 
        I121_un1_Y, N437, N436, N433, N432, N429, N327, N326, N333, 
        N329, N332, N335, \state_RNO_7[0] , \inf_abs1_a_1[2] , 
        \inf_abs0_a_0[2] , \state_RNO_8[1] , \inf_abs0_a_0[12] , N_3_0, 
        \DWACT_FINC_E[2] , \DWACT_FINC_E[5] , N_4, \DWACT_FINC_E[3] , 
        N_6, N_7, N_8, \DWACT_FINC_E[1] , N_9, N_11, N_3_1, 
        \DWACT_FINC_E_0[2] , \DWACT_FINC_E_0[5] , N_4_0, 
        \DWACT_FINC_E_0[3] , N_6_0, N_7_0, N_8_0, \DWACT_FINC_E_0[1] , 
        N_9_0, N_11_0, GND, VCC;
    
    OR2 un1_integ_0_0_ADD_26x26_fast_I56_Y (.A(I56_un1_Y), .B(N344), 
        .Y(N424));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I148_un1_Y (.A(N479), .B(N472), 
        .Y(I148_un1_Y));
    NOR2 inf_abs1_a_1_I_15 (.A(sr_old[4]), .B(sr_old[3]), .Y(
        \DWACT_FINC_E[1] ));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I58_un1_Y (.A(integral[7]), .B(
        \un1_next_int[7] ), .C(N342), .Y(I58_un1_Y));
    XNOR2 inf_abs1_a_1_I_23 (.A(sr_old[8]), .B(N_6), .Y(
        \inf_abs1_a_1[8] ));
    DFN1C0 \state[0]  (.D(\state_RNO_7[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[0]_net_1 ));
    XNOR2 inf_abs1_a_1_I_17 (.A(sr_old[6]), .B(N_8), .Y(
        \inf_abs1_a_1[6] ));
    DFN1E0C0 \integ[13]  (.D(\un1_integ[13] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[13]));
    NOR3C \state_RNIF0PH4[1]  (.A(sr_old[12]), .B(\state[1]_net_1 ), 
        .C(\inf_abs1_a_1[10] ), .Y(\inf_abs1_m[10] ));
    DFN1E0C0 \integ[24]  (.D(\un1_integ[24] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[24]));
    OR2 \state_RNII5U5A[0]  (.A(\un1_next_int_iv_1[11] ), .B(
        \un2_next_int_m[11] ), .Y(\un1_next_int[11] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I61_Y (.A(integral[7]), .B(
        \un1_next_int[7] ), .C(N336), .Y(N429));
    NOR3B inf_abs0_a_0_I_19 (.A(\DWACT_FINC_E_0[2] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[6]), .Y(N_7_0));
    OA1A \state_RNIO6755[1]  (.A(sr_old[12]), .B(\inf_abs1_a_1[12] ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[12] ));
    OR2 \state_RNI0HB66[0]  (.A(\un1_next_int_iv_1[4] ), .B(
        \inf_abs1_m[4] ), .Y(\un1_next_int[4] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I248_Y_0 (.A(integral[18]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I248_Y_0));
    NOR2A \state_RNI02011[1]  (.A(next_int_1_sqmuxa_1), .B(sr_old[3]), 
        .Y(\un18_next_int_m[3] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I172_un1_Y (.A(N467), .B(
        I144_un1_Y), .C(N506), .Y(I172_un1_Y));
    NOR3B inf_abs0_a_0_I_16 (.A(\DWACT_FINC_E_0[1] ), .B(
        \DWACT_FINC_E[0] ), .C(sr_new[5]), .Y(N_8_0));
    INV \integ_RNIH77A[24]  (.A(integral[24]), .Y(integral_i[24]));
    AO1B un1_integ_0_0_ADD_26x26_fast_I41_Y (.A(integral[17]), .B(
        integral[16]), .C(\un1_next_int_0_iv_0[13] ), .Y(N409));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I204_un1_Y (.A(N518), .B(N502), 
        .C(N655), .Y(I204_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I86_Y (.A(N408), .B(N404), .Y(
        N457));
    OR2 \state_RNIS3I11[1]  (.A(next_int_1_sqmuxa), .B(
        next_int_0_sqmuxa_1), .Y(\un1_next_int_0_iv_0[13] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I98_Y (.A(N420), .B(N417), .C(
        N416), .Y(N469));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I176_un1_Y (.A(N510), .B(N525), 
        .Y(I176_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I205_un1_Y_0 (.A(N466), .B(N474)
        , .C(N504), .Y(ADD_26x26_fast_I205_un1_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I150_un1_Y (.A(N481), .B(N474), 
        .Y(I150_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I51_Y (.A(N354), .B(N351), .Y(
        N419));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y (.A(
        ADD_26x26_fast_I230_Y_0), .B(\un1_next_int[0] ), .Y(
        \un1_integ[0] ));
    NOR2B inf_abs1_a_1_I_34 (.A(\DWACT_FINC_E_0[7] ), .B(
        \DWACT_FINC_E_0[6] ), .Y(N_2_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I144_un1_Y (.A(N419), .B(N415), 
        .C(N475), .Y(I144_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I253_Y (.A(I172_un1_Y), .B(
        ADD_26x26_fast_I206_Y_2), .C(ADD_26x26_fast_I253_Y_0), .Y(
        \un1_integ[23] ));
    DFN1E0C0 \integ[21]  (.D(\un1_integ[21] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[21]));
    XNOR2 inf_abs1_a_1_I_7 (.A(sr_old[2]), .B(N_12_0), .Y(
        \inf_abs1_a_1[2] ));
    DFN1E0C0 \integ_1[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral_1_0));
    OR3 un1_integ_0_0_ADD_26x26_fast_I205_Y (.A(I170_un1_Y), .B(
        ADD_26x26_fast_I205_Y_2), .C(I205_un1_Y), .Y(N619));
    OA1 un1_integ_0_0_ADD_26x26_fast_I190_un1_Y (.A(N487), .B(
        I162_un1_Y), .C(N526), .Y(I190_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I146_Y (.A(I146_un1_Y), .B(N469), 
        .Y(N523));
    NOR2B \state_RNI4KSN1[1]  (.A(\inf_abs1_a_1[2] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[2] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I142_Y (.A(I142_un1_Y), .B(N465), 
        .Y(N519));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I244_Y_0 (.A(integral[14]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I244_Y_0));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I231_Y (.A(
        ADD_26x26_fast_I231_Y_0), .B(N442), .Y(\un1_integ[1] ));
    AND3 inf_abs1_a_1_I_24 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E_0[4] ));
    XNOR2 inf_abs1_a_1_I_32 (.A(sr_old[11]), .B(N_3_0), .Y(
        \inf_abs1_a_1[11] ));
    DFN1E0C0 \integ[15]  (.D(\un1_integ[15] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[15]));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I213_un1_Y (.A(N466), .B(N474), 
        .C(ADD_26x26_fast_I213_un1_Y_0), .Y(I213_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I103_Y (.A(N348), .B(N351), .C(
        N425), .Y(N474));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I125_Y (.A(N399), .B(
        ADD_26x26_fast_I125_Y_0), .C(N456), .Y(N502));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_1 (.A(
        ADD_26x26_fast_I209_un1_Y_0), .B(N528), .C(
        ADD_26x26_fast_I209_Y_0), .Y(ADD_26x26_fast_I209_Y_1));
    AO1 un1_integ_0_0_ADD_26x26_fast_I94_Y (.A(N416), .B(N413), .C(
        N412), .Y(N465));
    NOR2 inf_abs0_a_0_I_6 (.A(sr_new[0]), .B(sr_new[1]), .Y(N_12));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I151_Y (.A(N474), .B(N482), .Y(
        N528));
    AND3 inf_abs1_a_1_I_22 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_6));
    OR2 un1_integ_0_0_ADD_26x26_fast_I74_Y (.A(I74_un1_Y), .B(N317), 
        .Y(N442));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I238_Y (.A(N658), .B(
        ADD_26x26_fast_I238_Y_0), .Y(\un1_integ[8] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I121_Y (.A(I121_un1_Y), .B(N440), 
        .Y(N493));
    NOR2B \state_RNIRTRQ3[1]  (.A(\inf_abs1[6]_net_1 ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[6] ));
    XA1 \state_RNI90H51[0]  (.A(sr_new[12]), .B(\inf_abs0[1]_net_1 ), 
        .C(\state[0]_net_1 ), .Y(\un1_next_int_iv_1[1] ));
    NOR3 inf_abs0_a_0_I_10 (.A(sr_new[0]), .B(sr_new[2]), .C(sr_new[1])
        , .Y(\DWACT_FINC_E[0] ));
    NOR2A \state_RNIRLHL_0[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), 
        .Y(next_int_1_sqmuxa_1));
    OR3 un1_integ_0_0_ADD_26x26_fast_I5_P0N (.A(\un2_next_int_m[5] ), 
        .B(\un1_next_int_iv_1[5] ), .C(\integ[5]_net_1 ), .Y(N333));
    NOR2A \state_RNI57011[1]  (.A(next_int_1_sqmuxa_1), .B(sr_old[8]), 
        .Y(\un18_next_int_m[8] ));
    NOR2A \state_RNI1E0C[0]  (.A(\state[0]_net_1 ), .B(sr_new[12]), .Y(
        next_int_1_sqmuxa));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I246_Y (.A(
        \un1_next_int_0_iv[13] ), .B(integral[16]), .C(N635), .Y(
        \un1_integ[16] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I252_Y_0 (.A(integral[22]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I252_Y_0));
    NOR2B \state_RNIRLHL[1]  (.A(\state[1]_net_1 ), .B(sr_old[12]), .Y(
        next_int_0_sqmuxa_1));
    NOR2B \state_RNIG1PH4[1]  (.A(\inf_abs1[8]_net_1 ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[8] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I39_Y (.A(integral[17]), .B(
        integral[18]), .C(\un1_next_int_0_iv_0[13] ), .Y(N407));
    OA1B un1_integ_0_0_ADD_26x26_fast_I32_Y (.A(integral[21]), .B(
        integral[20]), .C(\un1_next_int_0_iv_0[13] ), .Y(N400));
    OR3 un1_integ_0_0_ADD_26x26_fast_I213_Y (.A(I186_un1_Y), .B(N519), 
        .C(I213_un1_Y), .Y(N635));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I194_un1_Y (.A(N534), .B(N442), 
        .Y(I194_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I108_un1_Y (.A(N430), .B(N427), 
        .Y(I108_un1_Y));
    NOR2A inf_abs0_a_0_I_11 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .Y(
        N_10));
    AO1B un1_integ_0_0_ADD_26x26_fast_I125_Y_0 (.A(integral[23]), .B(
        integral[24]), .C(\un1_next_int_0_iv_0[13] ), .Y(
        ADD_26x26_fast_I125_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I211_Y_1_0 (.A(N462), .B(N470), 
        .Y(ADD_26x26_fast_I211_Y_1_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I100_Y (.A(N422), .B(N419), .C(
        N418), .Y(N471));
    OR3 un1_integ_0_0_ADD_26x26_fast_I12_P0N (.A(\un2_next_int_m[12] ), 
        .B(\un1_next_int_iv_0[12] ), .C(integral[12]), .Y(N354));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I10_G0N (.A(\un1_next_int[10] ), 
        .B(integral[10]), .Y(N347));
    DFN1E0C0 \integ[12]  (.D(\un1_integ[12] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[12]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I109_Y (.A(N431), .B(N427), .Y(
        N480));
    AO1A \state_RNI1NU44[1]  (.A(\inf_abs1[2]_net_1 ), .B(
        next_int_1_sqmuxa_1), .C(\inf_abs1_m[2] ), .Y(
        \un1_next_int_iv_0[2] ));
    XNOR2 inf_abs1_a_1_I_35 (.A(sr_old[12]), .B(N_2_0), .Y(
        \inf_abs1_a_1[12] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I205_Y_0 (.A(integral[23]), .B(
        integral[22]), .C(\un1_next_int_0_iv_0[13] ), .Y(
        ADD_26x26_fast_I205_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I115_Y (.A(N433), .B(N437), .Y(
        N486));
    OA1 un1_integ_0_0_ADD_26x26_fast_I12_G0N (.A(\un2_next_int_m[12] ), 
        .B(\un1_next_int_iv_0[12] ), .C(integral[12]), .Y(N353));
    OR2 un1_integ_0_0_ADD_26x26_fast_I208_Y_0 (.A(N455), .B(N463), .Y(
        ADD_26x26_fast_I208_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I111_Y (.A(N429), .B(N433), .Y(
        N482));
    NOR2A inf_abs1_a_1_I_25 (.A(\DWACT_FINC_E_0[4] ), .B(sr_old[8]), 
        .Y(N_5_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I2_P0N (.A(\un1_next_int[2] ), .B(
        \integ[2]_net_1 ), .Y(N324));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I250_Y_0 (.A(integral[20]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I250_Y_0));
    NOR3A inf_abs1_a_1_I_27 (.A(\DWACT_FINC_E_0[4] ), .B(sr_old[8]), 
        .C(sr_old[9]), .Y(N_4));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I142_un1_Y (.A(N473), .B(N466), 
        .Y(I142_un1_Y));
    NOR3B \state_RNI71AB2[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[10]_net_1 ), .Y(\un2_next_int_m[10] ));
    DFN1E0C0 \integ[10]  (.D(\un1_integ[10] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[10]));
    OA1 un1_integ_0_0_ADD_26x26_fast_I188_un1_Y (.A(N483), .B(
        I160_un1_Y), .C(N522), .Y(I188_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I180_un1_Y (.A(N514), .B(N529), 
        .Y(I180_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I6_G0N (.A(\un1_next_int[6] ), 
        .B(integral[6]), .Y(N335));
    NOR2B \state_RNI06J52_0[0]  (.A(\inf_abs0[7]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[7] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I249_Y (.A(I210_un1_Y), .B(
        ADD_26x26_fast_I210_Y_1), .C(ADD_26x26_fast_I249_Y_0), .Y(
        \un1_integ[19] ));
    GND GND_i (.Y(GND));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I146_un1_Y (.A(N477), .B(N470), 
        .Y(I146_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I6_P0N (.A(\un1_next_int[6] ), .B(
        integral[6]), .Y(N336));
    NOR2A \state_RNI35011[1]  (.A(next_int_1_sqmuxa_1), .B(sr_old[6]), 
        .Y(\un18_next_int_m[6] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I1_G0N (.A(\un1_next_int_iv_0[1] )
        , .B(\un1_next_int_iv_1[1] ), .C(\integ[1]_net_1 ), .Y(N320));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I107_Y (.A(N429), .B(N425), .Y(
        N478));
    OR3 \state_RNID1FE3[0]  (.A(\inf_abs0_m[8] ), .B(
        \un18_next_int_m[8] ), .C(\un2_next_int_m[8] ), .Y(
        \un1_next_int_iv_1[8] ));
    NOR2B \state_RNIAUU33[1]  (.A(\inf_abs1[4]_net_1 ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[4] ));
    XNOR2 inf_abs1_a_1_I_9 (.A(sr_old[3]), .B(N_11), .Y(
        \inf_abs1_a_1[3] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I38_Y (.A(integral[17]), .B(
        integral[18]), .C(\un1_next_int_0_iv_0[13] ), .Y(N406));
    OA1 un1_integ_0_0_ADD_26x26_fast_I209_un1_Y_0 (.A(N489), .B(
        I163_un1_Y), .C(N512), .Y(ADD_26x26_fast_I209_un1_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I255_Y (.A(I204_un1_Y), .B(
        ADD_26x26_fast_I204_Y_3), .C(ADD_26x26_fast_I255_Y_0), .Y(
        \un1_integ[25] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I204_Y_0 (.A(integral[24]), .B(
        integral[23]), .C(\un1_next_int_0_iv[13] ), .Y(
        ADD_26x26_fast_I204_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I243_Y (.A(N525), .B(I190_un1_Y), 
        .C(ADD_26x26_fast_I243_Y_0), .Y(\un1_integ[13] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I231_Y_0 (.A(
        \un1_next_int_iv_0[1] ), .B(\un1_next_int_iv_1[1] ), .C(
        \integ[1]_net_1 ), .Y(ADD_26x26_fast_I231_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I69_Y (.A(N324), .B(N327), .Y(
        N437));
    AO1 un1_integ_0_0_ADD_26x26_fast_I62_Y (.A(N332), .B(N336), .C(
        N335), .Y(N430));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I193_un1_Y (.A(N478), .B(N486), 
        .C(N493), .Y(I193_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I153_Y (.A(N484), .B(N476), .Y(
        N530));
    XA1A \state_RNIOMJ12[1]  (.A(sr_old[12]), .B(\inf_abs1[1]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[1] ));
    XNOR2 inf_abs0_a_0_I_7 (.A(sr_new[2]), .B(N_12), .Y(
        \inf_abs0_a_0[2] ));
    OA1A un1_integ_0_0_ADD_26x26_fast_I49_Y (.A(
        \un1_next_int_0_iv[13] ), .B(integral[13]), .C(N354), .Y(N417));
    OA1B un1_integ_0_0_ADD_26x26_fast_I42_Y (.A(integral[15]), .B(
        integral[16]), .C(\un1_next_int_0_iv_0[13] ), .Y(N410));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I145_Y (.A(N419), .B(N415), .C(
        N476), .Y(N522));
    MX2 \inf_abs1[4]  (.A(sr_old[4]), .B(\inf_abs1_a_1[4] ), .S(
        sr_old[12]), .Y(\inf_abs1[4]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I10_P0N (.A(\un1_next_int[10] ), 
        .B(integral[10]), .Y(N348));
    NOR2B \state_RNIJIBH[0]  (.A(sr_new[9]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[9] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I1_P0N (.A(\un1_next_int_iv_0[1] )
        , .B(\un1_next_int_iv_1[1] ), .C(\integ[1]_net_1 ), .Y(N321));
    OA1 un1_integ_0_0_ADD_26x26_fast_I184_un1_Y (.A(N479), .B(
        I156_un1_Y), .C(N518), .Y(I184_un1_Y));
    NOR3B \state_RNIM83S1[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[8] ), .Y(\un2_next_int_m[8] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I192_un1_Y (.A(N530), .B(N491), 
        .Y(I192_un1_Y));
    NOR3A inf_abs0_a_0_I_13 (.A(\DWACT_FINC_E[0] ), .B(sr_new[3]), .C(
        sr_new[4]), .Y(N_9_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I156_un1_Y (.A(N487), .B(N480), 
        .Y(I156_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I141_Y (.A(N464), .B(N472), .Y(
        N518));
    NOR2B \state_RNI3UFB2_0[0]  (.A(\inf_abs0[11]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[11] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I93_Y (.A(N411), .B(N415), .Y(
        N464));
    AO1B un1_integ_0_0_ADD_26x26_fast_I37_Y (.A(integral[18]), .B(
        integral[19]), .C(\un1_next_int_0_iv_0[13] ), .Y(N405));
    OR3 un1_integ_0_0_ADD_26x26_fast_I194_Y (.A(N479), .B(I156_un1_Y), 
        .C(I194_un1_Y), .Y(N655));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I0_G0N (.A(N_3), .B(
        \integ[0]_net_1 ), .Y(N317));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I73_Y (.A(N318), .B(N321), .Y(
        N441));
    OA1 un1_integ_0_0_ADD_26x26_fast_I59_Y (.A(integral[7]), .B(
        \un1_next_int[7] ), .C(N342), .Y(N427));
    AO1 un1_integ_0_0_ADD_26x26_fast_I52_Y (.A(N347), .B(N351), .C(
        N350), .Y(N420));
    NOR2A \state_RNO[1]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 ), 
        .Y(\state_RNO_8[1] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I34_Y (.A(integral[20]), .B(
        integral[19]), .C(\un1_next_int_0_iv_0[13] ), .Y(N402));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I236_Y (.A(\un1_next_int[6] ), 
        .B(integral[6]), .C(N539), .Y(\un1_integ[6] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I54_un1_Y (.A(N344), .B(N348), 
        .Y(I54_un1_Y));
    OR2 \state_RNIF7EQ7[1]  (.A(\un1_next_int_iv_0[11] ), .B(
        \inf_abs0_m[11] ), .Y(\un1_next_int_iv_1[11] ));
    NOR2A \state_RNI68011[1]  (.A(next_int_1_sqmuxa_1), .B(sr_old[9]), 
        .Y(\un18_next_int_m[9] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I150_Y (.A(I150_un1_Y), .B(N473), 
        .Y(N527));
    DFN1E0C0 \integ[0]  (.D(\un1_integ[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(\integ[0]_net_1 ));
    OR2 \state_RNINV523[1]  (.A(\un1_next_int_iv_1[0] ), .B(
        \un1_next_int_iv_0[0] ), .Y(\un1_next_int[0] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I120_Y (.A(I120_un1_Y), .B(N438), 
        .Y(N491));
    AO1 un1_integ_0_0_ADD_26x26_fast_I104_Y (.A(N426), .B(N423), .C(
        N422), .Y(N475));
    VCC VCC_i (.Y(VCC));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I129_Y (.A(N403), .B(N399), .C(
        N460), .Y(N506));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I113_Y (.A(N431), .B(N435), .Y(
        N484));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I241_Y_0 (.A(\un1_next_int[11] ), 
        .B(integral[11]), .Y(ADD_26x26_fast_I241_Y_0));
    XNOR2 inf_abs0_a_0_I_28 (.A(sr_new[10]), .B(N_4_0), .Y(
        \inf_abs0_a_0[10] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I89_Y (.A(N411), .B(N407), .Y(
        N460));
    AO1 un1_integ_0_0_ADD_26x26_fast_I68_Y (.A(N323), .B(N327), .C(
        N326), .Y(N436));
    AO1 un1_integ_0_0_ADD_26x26_fast_I211_Y_0 (.A(N469), .B(N462), .C(
        N461), .Y(ADD_26x26_fast_I211_Y_0));
    DFN1E0C0 \integ[4]  (.D(\un1_integ[4] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(\integ[4]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I108_Y (.A(I108_un1_Y), .B(N426), 
        .Y(N479));
    NOR2 \state_RNIB3LN_0[1]  (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(N_46_1_0));
    NOR3 inf_abs1_a_1_I_18 (.A(sr_old[5]), .B(sr_old[4]), .C(sr_old[3])
        , .Y(\DWACT_FINC_E[2] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I3_G0N (.A(\un1_next_int_iv_0[3] )
        , .B(\un1_next_int_iv_1[3] ), .C(\integ[3]_net_1 ), .Y(N326));
    AO13 un1_integ_0_0_ADD_26x26_fast_I48_Y (.A(integral[13]), .B(N353)
        , .C(\un1_next_int_0_iv[13] ), .Y(N416));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I195_un1_Y (.A(N482), .B(N490), 
        .C(\un1_next_int[0] ), .Y(I195_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I102_un1_Y (.A(N348), .B(N351), 
        .C(N424), .Y(I102_un1_Y));
    DFN1E0C0 \integ[3]  (.D(\un1_integ[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(\integ[3]_net_1 ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I252_Y (.A(I174_un1_Y), .B(
        ADD_26x26_fast_I207_Y_2), .C(ADD_26x26_fast_I252_Y_0), .Y(
        \un1_integ[22] ));
    DFN1E0C0 \integ[6]  (.D(\un1_integ[6] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(integral[6]));
    XNOR2 inf_abs0_a_0_I_14 (.A(sr_new[5]), .B(N_9_0), .Y(
        \inf_abs0_a_0[5] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I210_Y_1 (.A(I136_un1_Y), .B(N459)
        , .C(I180_un1_Y), .Y(ADD_26x26_fast_I210_Y_1));
    AND3 inf_abs0_a_0_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[5] ), .Y(
        \DWACT_FINC_E[6] ));
    NOR2A \state_RNI24011[1]  (.A(next_int_1_sqmuxa_1), .B(sr_old[5]), 
        .Y(\un18_next_int_m[5] ));
    XOR3 un1_integ_0_0_ADD_26x26_fast_I239_Y (.A(\un1_next_int[9] ), 
        .B(integral[9]), .C(N655), .Y(\un1_integ[9] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I106_un1_Y (.A(N428), .B(N425), 
        .Y(I106_un1_Y));
    OR2 \state_RNIMIC23[0]  (.A(\un1_next_int_iv_0[4] ), .B(
        \un2_next_int_m[4] ), .Y(\un1_next_int_iv_1[4] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I58_Y (.A(\un1_next_int[8] ), .B(
        integral[8]), .C(I58_un1_Y), .Y(N426));
    NOR3B \state_RNI721G1[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[4] ), .Y(\un2_next_int_m[4] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I67_Y (.A(\integ[4]_net_1 ), .B(
        \un1_next_int[4] ), .C(N327), .Y(N435));
    XNOR2 inf_abs0_a_0_I_12 (.A(sr_new[4]), .B(N_10), .Y(
        \inf_abs0_a_0[4] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I253_Y_0 (.A(integral[23]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I253_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I157_Y (.A(N488), .B(N480), .Y(
        N534));
    AO1 un1_integ_0_0_ADD_26x26_fast_I64_Y (.A(N329), .B(N333), .C(
        N332), .Y(N432));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I50_un1_Y (.A(N350), .B(N354), 
        .Y(I50_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I212_un1_Y (.A(N534), .B(N442), 
        .C(N518), .Y(I212_un1_Y));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I127_Y (.A(N401), .B(
        ADD_26x26_fast_I127_Y_0), .C(N458), .Y(N504));
    AO1 un1_integ_0_0_ADD_26x26_fast_I110_Y (.A(N432), .B(N429), .C(
        N428), .Y(N481));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I211_un1_Y_0 (.A(N478), .B(N486)
        , .C(N493), .Y(ADD_26x26_fast_I211_un1_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I90_Y (.A(N408), .B(N412), .Y(
        N461));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I233_Y (.A(
        ADD_26x26_fast_I233_Y_0), .B(N491), .Y(\un1_integ[3] ));
    NOR3A inf_abs0_a_0_I_31 (.A(\DWACT_FINC_E[6] ), .B(sr_new[9]), .C(
        sr_new[10]), .Y(N_3_1));
    AO1B un1_integ_0_0_ADD_26x26_fast_I47_Y (.A(integral[13]), .B(
        integral[14]), .C(\un1_next_int_0_iv[13] ), .Y(N415));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I119_Y (.A(N441), .B(N437), .Y(
        N490));
    MX2 \inf_abs0[7]  (.A(sr_new[7]), .B(\inf_abs0_a_0[7] ), .S(
        sr_new_0_0), .Y(\inf_abs0[7]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I70_Y (.A(N320), .B(N324), .C(
        N323), .Y(N438));
    DFN1E0C0 \integ[5]  (.D(\un1_integ[5] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(\integ[5]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I161_Y (.A(N486), .B(N493), .C(
        N485), .Y(N539));
    OA1B un1_integ_0_0_ADD_26x26_fast_I44_Y (.A(integral[14]), .B(
        integral[15]), .C(\un1_next_int_0_iv_0[13] ), .Y(N412));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I245_Y (.A(
        \un1_next_int_0_iv[13] ), .B(integral[15]), .C(N637), .Y(
        \un1_integ[15] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I95_Y (.A(N413), .B(N417), .Y(
        N466));
    DFN1E0C0 \integ[2]  (.D(\un1_integ[2] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(\integ[2]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I135_Y (.A(N458), .B(N466), .Y(
        N512));
    OR2 un1_integ_0_0_ADD_26x26_fast_I88_Y (.A(N410), .B(N406), .Y(
        N459));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I247_Y (.A(
        \un1_next_int_0_iv[13] ), .B(integral[17]), .C(N633), .Y(
        \un1_integ[17] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I237_Y_0 (.A(integral[7]), .B(
        \un1_next_int[7] ), .Y(ADD_26x26_fast_I237_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I57_Y (.A(N342), .B(N345), .Y(
        N425));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I186_un1_Y (.A(N466), .B(N474), 
        .C(N535), .Y(I186_un1_Y));
    NOR3 inf_abs0_a_0_I_29 (.A(sr_new[7]), .B(sr_new[6]), .C(sr_new[8])
        , .Y(\DWACT_FINC_E_0[5] ));
    DFN1E0C0 \integ[23]  (.D(\un1_integ[23] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[23]));
    OR2 un1_integ_0_0_ADD_26x26_fast_I8_P0N (.A(\un1_next_int[8] ), .B(
        integral[8]), .Y(N342));
    OR3 un1_integ_0_0_ADD_26x26_fast_I212_Y (.A(I184_un1_Y), .B(N517), 
        .C(I212_un1_Y), .Y(N633));
    AO1 un1_integ_0_0_ADD_26x26_fast_I206_Y_2 (.A(
        ADD_26x26_fast_I206_un1_Y_0), .B(N522), .C(
        ADD_26x26_fast_I206_Y_1), .Y(ADD_26x26_fast_I206_Y_2));
    OR2 un1_integ_0_0_ADD_26x26_fast_I54_Y (.A(I54_un1_Y), .B(N347), 
        .Y(N422));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I131_Y (.A(N401), .B(N405), .C(
        N462), .Y(N508));
    XNOR2 inf_abs0_a_0_I_26 (.A(sr_new[9]), .B(N_5), .Y(
        \inf_abs0_a_0[9] ));
    NOR3B inf_abs1_a_1_I_19 (.A(\DWACT_FINC_E[2] ), .B(
        \DWACT_FINC_E_0[0] ), .C(sr_old[6]), .Y(N_7));
    NOR3B \state_RNI3UFB2[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[11]_net_1 ), .Y(\un2_next_int_m[11] ));
    NOR3B inf_abs1_a_1_I_16 (.A(\DWACT_FINC_E[1] ), .B(
        \DWACT_FINC_E_0[0] ), .C(sr_old[5]), .Y(N_8));
    XNOR3 un1_integ_0_0_ADD_26x26_fast_I254_Y (.A(
        \un1_next_int_0_iv[13] ), .B(integral[24]), .C(N619), .Y(
        \un1_integ[24] ));
    DFN1E0C0 \integ[19]  (.D(\un1_integ[19] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[19]));
    NOR2 inf_abs0_a_0_I_15 (.A(sr_new[3]), .B(sr_new[4]), .Y(
        \DWACT_FINC_E_0[1] ));
    NOR2A \state_RNI13011[1]  (.A(next_int_1_sqmuxa_1), .B(sr_old[4]), 
        .Y(\un18_next_int_m[4] ));
    MX2 \inf_abs1[8]  (.A(sr_old[8]), .B(\inf_abs1_a_1[8] ), .S(
        sr_old[12]), .Y(\inf_abs1[8]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I117_Y (.A(N439), .B(N435), .Y(
        N488));
    DFN1E0C0 \integ[17]  (.D(\un1_integ[17] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[17]));
    XOR2 inf_abs0_a_0_I_5 (.A(sr_new[0]), .B(sr_new[1]), .Y(
        \inf_abs0_a_0[1] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I33_Y (.A(integral[21]), .B(
        integral[20]), .C(\un1_next_int_0_iv_0[13] ), .Y(N401));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I255_Y_0 (.A(integral[25]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I255_Y_0));
    AO1B un1_integ_0_0_ADD_26x26_fast_I127_Y_0 (.A(integral[22]), .B(
        integral[23]), .C(\un1_next_int_0_iv[13] ), .Y(
        ADD_26x26_fast_I127_Y_0));
    NOR2B \state_RNIEDBH[0]  (.A(sr_new[4]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[4] ));
    DFN1E0C0 \integ[14]  (.D(\un1_integ[14] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[14]));
    XNOR2 inf_abs0_a_0_I_17 (.A(sr_new[6]), .B(N_8_0), .Y(
        \inf_abs0_a_0[6] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I87_Y (.A(N409), .B(N405), .Y(
        N458));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y_0 (.A(\integ[2]_net_1 ), 
        .B(\un1_next_int[2] ), .Y(ADD_26x26_fast_I232_Y_0));
    MX2 \inf_abs1[0]  (.A(sr_old[0]), .B(sr_old[0]), .S(sr_old[12]), 
        .Y(\inf_abs1[0]_net_1 ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I84_Y (.A(N406), .B(N402), .Y(
        N455));
    AO1 un1_integ_0_0_ADD_26x26_fast_I154_Y (.A(N485), .B(N478), .C(
        N477), .Y(N531));
    MX2 \inf_abs1[11]  (.A(sr_old[11]), .B(\inf_abs1_a_1[11] ), .S(
        sr_old[12]), .Y(\inf_abs1[11]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I11_G0N (.A(\un1_next_int[11] ), 
        .B(integral[11]), .Y(N350));
    MX2 \inf_abs1[2]  (.A(sr_old[2]), .B(\inf_abs1_a_1[2] ), .S(
        sr_old[12]), .Y(\inf_abs1[2]_net_1 ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I140_Y (.A(N471), .B(N464), .C(
        N463), .Y(N517));
    NOR2B \state_RNIMR7Q2[1]  (.A(\inf_abs1_a_1[5] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[5] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I149_Y (.A(N480), .B(N472), .Y(
        N526));
    AO1 un1_integ_0_0_ADD_26x26_fast_I158_Y (.A(N489), .B(N482), .C(
        N481), .Y(N535));
    NOR3B \state_RNI8DE12[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[9] ), .Y(\un2_next_int_m[9] ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I249_Y_0 (.A(integral[19]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I249_Y_0));
    DFN1E0C0 \integ[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[25]));
    NOR3B \state_RNIQ2MA1[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[3] ), .Y(\un2_next_int_m[3] ));
    NOR3B \state_RNIPALQ[0]  (.A(\state[0]_net_1 ), .B(sr_new_0_0), .C(
        sr_new[0]), .Y(\un2_next_int_m[0] ));
    MX2 \inf_abs1[6]  (.A(sr_old[6]), .B(\inf_abs1_a_1[6] ), .S(
        sr_old[12]), .Y(\inf_abs1[6]_net_1 ));
    NOR3 inf_abs0_a_0_I_33 (.A(sr_new[10]), .B(sr_new[9]), .C(
        sr_new[11]), .Y(\DWACT_FINC_E[7] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I230_Y_0 (.A(\integ[0]_net_1 ), 
        .B(N_3), .Y(ADD_26x26_fast_I230_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I242_Y (.A(N527), .B(I191_un1_Y), 
        .C(ADD_26x26_fast_I242_Y_0), .Y(\un1_integ[12] ));
    XNOR2 inf_abs0_a_0_I_20 (.A(sr_new[7]), .B(N_7_0), .Y(
        \inf_abs0_a_0[7] ));
    DFN1E0C0 \integ[11]  (.D(\un1_integ[11] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1_0), .Q(integral[11]));
    DFN1E0C0 \integ[16]  (.D(\un1_integ[16] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[16]));
    XNOR2 inf_abs1_a_1_I_28 (.A(sr_old[10]), .B(N_4), .Y(
        \inf_abs1_a_1[10] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I211_Y_1 (.A(
        ADD_26x26_fast_I211_un1_Y_0), .B(N531), .C(
        ADD_26x26_fast_I211_Y_1_0), .Y(ADD_26x26_fast_I211_Y_1));
    NOR3 inf_abs1_a_1_I_10 (.A(sr_old[1]), .B(sr_old[0]), .C(sr_old[2])
        , .Y(\DWACT_FINC_E_0[0] ));
    OR2 \state_RNIBQL7A[0]  (.A(\un1_next_int_iv_1[10] ), .B(
        \un2_next_int_m[10] ), .Y(\un1_next_int[10] ));
    MX2B un1_next_int_0_sqmuxa_0__m2 (.A(sr_new_0_0), .B(sr_old[12]), 
        .S(\state[1]_net_1 ), .Y(N_3));
    OR2 un1_integ_0_0_ADD_26x26_fast_I96_Y (.A(I96_un1_Y), .B(N414), 
        .Y(N467));
    MX2 \inf_abs0[10]  (.A(sr_new[10]), .B(\inf_abs0_a_0[10] ), .S(
        sr_new_0_0), .Y(\inf_abs0[10]_net_1 ));
    OR2 \state_RNIJKBI1[0]  (.A(\un18_next_int_m[6] ), .B(
        \inf_abs0_m[6] ), .Y(\un1_next_int_iv_0[6] ));
    NOR2B \state_RNIGFBH[0]  (.A(sr_new[6]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[6] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I2_G0N (.A(\un1_next_int[2] ), 
        .B(\integ[2]_net_1 ), .Y(N323));
    NOR2B \state_RNISU184[1]  (.A(\inf_abs1_a_1[9] ), .B(
        next_int_0_sqmuxa_1), .Y(\inf_abs1_m[9] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I114_Y (.A(N436), .B(N433), .C(
        N432), .Y(N485));
    OR2 \state_RNIT2808[0]  (.A(\un1_next_int_iv_1[8] ), .B(
        \inf_abs1_m[8] ), .Y(\un1_next_int[8] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I189_un1_Y (.A(N524), .B(N539), 
        .Y(I189_un1_Y));
    MX2 \inf_abs1[1]  (.A(sr_old[1]), .B(\inf_abs1_a_1[1] ), .S(
        sr_old[12]), .Y(\inf_abs1[1]_net_1 ));
    NOR2 inf_abs0_a_0_I_21 (.A(sr_new[6]), .B(sr_new[7]), .Y(
        \DWACT_FINC_E_0[3] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I147_Y (.A(N478), .B(N470), .Y(
        N524));
    DFN1E0C0 \integ[9]  (.D(\un1_integ[9] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(integral[9]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I242_Y_0 (.A(
        \un2_next_int_m[12] ), .B(\un1_next_int_iv_0[12] ), .C(
        integral[12]), .Y(ADD_26x26_fast_I242_Y_0));
    AX1D un1_integ_0_0_ADD_26x26_fast_I235_Y (.A(N487), .B(I162_un1_Y), 
        .C(ADD_26x26_fast_I235_Y_0), .Y(\un1_integ[5] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I63_Y (.A(N333), .B(N336), .Y(
        N431));
    NOR2A inf_abs1_a_1_I_11 (.A(\DWACT_FINC_E_0[0] ), .B(sr_old[3]), 
        .Y(N_10_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I96_un1_Y (.A(N418), .B(N415), 
        .Y(I96_un1_Y));
    AO1 un1_integ_0_0_ADD_26x26_fast_I118_Y (.A(N440), .B(N437), .C(
        N436), .Y(N489));
    AX1D un1_integ_0_0_ADD_26x26_fast_I237_Y (.A(N483), .B(I160_un1_Y), 
        .C(ADD_26x26_fast_I237_Y_0), .Y(\un1_integ[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I133_Y (.A(N464), .B(N456), .Y(
        N510));
    MX2 \inf_abs0[2]  (.A(sr_new[2]), .B(\inf_abs0_a_0[2] ), .S(
        sr_new_0_0), .Y(\inf_abs0[2]_net_1 ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I30_Y (.A(integral[22]), .B(
        integral[21]), .C(\un1_next_int_0_iv_0[13] ), .Y(N398));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I160_un1_Y (.A(N484), .B(N491), 
        .Y(I160_un1_Y));
    AO1 \state_RNI3K0C1[0]  (.A(sr_new[0]), .B(next_int_1_sqmuxa), .C(
        \un2_next_int_m[0] ), .Y(\un1_next_int_iv_1[0] ));
    DFN1E0C0 \integ[22]  (.D(\un1_integ[22] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[22]));
    NOR3 inf_abs1_a_1_I_8 (.A(sr_old[1]), .B(sr_old[0]), .C(sr_old[2]), 
        .Y(N_11));
    AO1B un1_integ_0_0_ADD_26x26_fast_I43_Y (.A(integral[16]), .B(
        integral[15]), .C(\un1_next_int_0_iv_0[13] ), .Y(N411));
    INV \integ_RNII87A[25]  (.A(integral[25]), .Y(integral_i[25]));
    DFN1E0C0 \integ_0[25]  (.D(\un1_integ[25] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral_0_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I192_Y (.A(N529), .B(I192_un1_Y), 
        .Y(N649));
    DFN1E0C0 \integ[1]  (.D(\un1_integ[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(\integ[1]_net_1 ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I35_Y (.A(integral[19]), .B(
        integral[20]), .C(\un1_next_int_0_iv_0[13] ), .Y(N403));
    NOR2B inf_abs0_a_0_I_34 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_2));
    NOR3B \state_RNI44NQ1[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[6] ), .Y(\un2_next_int_m[6] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I91_Y (.A(N409), .B(N413), .Y(
        N462));
    AX1D un1_integ_0_0_ADD_26x26_fast_I250_Y (.A(I178_un1_Y), .B(
        ADD_26x26_fast_I209_Y_1), .C(ADD_26x26_fast_I250_Y_0), .Y(
        \un1_integ[20] ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I240_Y_0 (.A(integral[10]), .B(
        \un1_next_int[10] ), .Y(ADD_26x26_fast_I240_Y_0));
    NOR2A \state_RNIEN8V[1]  (.A(next_int_1_sqmuxa_1), .B(sr_old[10]), 
        .Y(\un18_next_int_m[10] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I71_Y (.A(N324), .B(N321), .Y(
        N439));
    XA1A \state_RNI5FA64[1]  (.A(sr_old[12]), .B(\inf_abs1[7]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[7] ));
    DFN1E0C0 \integ[20]  (.D(\un1_integ[20] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[20]));
    AX1D un1_integ_0_0_ADD_26x26_fast_I244_Y (.A(N523), .B(I189_un1_Y), 
        .C(ADD_26x26_fast_I244_Y_0), .Y(\un1_integ[14] ));
    NOR3 inf_abs1_a_1_I_29 (.A(sr_old[7]), .B(sr_old[6]), .C(sr_old[8])
        , .Y(\DWACT_FINC_E[5] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I207_Y_1 (.A(N404), .B(N400), .C(
        N461), .Y(ADD_26x26_fast_I207_Y_1));
    OR2 un1_integ_0_0_ADD_26x26_fast_I106_Y (.A(I106_un1_Y), .B(N424), 
        .Y(N477));
    XNOR2 inf_abs0_a_0_I_32 (.A(sr_new[11]), .B(N_3_1), .Y(
        \inf_abs0_a_0[11] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I208_Y_1 (.A(
        ADD_26x26_fast_I208_un1_Y_0), .B(N526), .C(
        ADD_26x26_fast_I208_Y_0), .Y(ADD_26x26_fast_I208_Y_1));
    OR2 un1_integ_0_0_ADD_26x26_fast_I102_Y (.A(I102_un1_Y), .B(N420), 
        .Y(N473));
    AX1D un1_integ_0_0_ADD_26x26_fast_I251_Y (.A(I176_un1_Y), .B(
        ADD_26x26_fast_I208_Y_1), .C(ADD_26x26_fast_I251_Y_0), .Y(
        \un1_integ[21] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I121_un1_Y (.A(N441), .B(
        \un1_next_int[0] ), .Y(I121_un1_Y));
    XNOR2 inf_abs1_a_1_I_26 (.A(sr_old[9]), .B(N_5_0), .Y(
        \inf_abs1_a_1[9] ));
    DFN1E0C0 \integ[18]  (.D(\un1_integ[18] ), .CLK(clk_c), .CLR(
        n_rst_c), .E(N_46_1), .Q(integral[18]));
    NOR2B \state_RNIFEBH[0]  (.A(sr_new[5]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[5] ));
    OR3 \state_RNILPDQ5[0]  (.A(\inf_abs0_m[9] ), .B(
        \un18_next_int_m[9] ), .C(\inf_abs1_m[9] ), .Y(
        \un1_next_int_iv_1[9] ));
    OR3 \state_RNI7EJC4[0]  (.A(\inf_abs0_m[5] ), .B(
        \un18_next_int_m[5] ), .C(\inf_abs1_m[5] ), .Y(
        \un1_next_int_iv_1[5] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I209_Y_0 (.A(N465), .B(N458), .C(
        N457), .Y(ADD_26x26_fast_I209_Y_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I148_Y (.A(I148_un1_Y), .B(N471), 
        .Y(N525));
    XA1 \state_RNILURA1[0]  (.A(sr_new[12]), .B(\inf_abs0[2]_net_1 ), 
        .C(\state[0]_net_1 ), .Y(\un1_next_int_iv_1[2] ));
    NOR3B \state_RNIL2CL1[0]  (.A(sr_new_0_0), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[5] ), .Y(\un2_next_int_m[5] ));
    XA1A \state_RNIC9UE5[1]  (.A(sr_old[12]), .B(\inf_abs1[11]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[11] ));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I60_Y (.A(N335), .B(integral[7]), 
        .C(\un1_next_int[7] ), .Y(N428));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I232_Y (.A(
        ADD_26x26_fast_I232_Y_0), .B(N493), .Y(\un1_integ[2] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I204_Y_2 (.A(N398), .B(
        ADD_26x26_fast_I204_Y_0), .C(N455), .Y(ADD_26x26_fast_I204_Y_2)
        );
    DFN1C0 \state[1]  (.D(\state_RNO_8[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\state[1]_net_1 ));
    XNOR2 inf_abs0_a_0_I_23 (.A(sr_new[8]), .B(N_6_0), .Y(
        \inf_abs0_a_0[8] ));
    NOR2B \state_RNI71AB2_0[0]  (.A(\inf_abs0[10]_net_1 ), .B(
        next_int_1_sqmuxa), .Y(\inf_abs0_m[10] ));
    NOR3A inf_abs1_a_1_I_13 (.A(\DWACT_FINC_E_0[0] ), .B(sr_old[4]), 
        .C(sr_old[3]), .Y(N_9));
    MX2 \inf_abs1[7]  (.A(sr_old[7]), .B(\inf_abs1_a_1[7] ), .S(
        sr_old[12]), .Y(\inf_abs1[7]_net_1 ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I9_G0N (.A(\un1_next_int[9] ), 
        .B(integral[9]), .Y(N344));
    OA1B un1_integ_0_0_ADD_26x26_fast_I40_Y (.A(integral[16]), .B(
        integral[17]), .C(\un1_next_int_0_iv_0[13] ), .Y(N408));
    OA1 un1_integ_0_0_ADD_26x26_fast_I65_Y (.A(\integ[4]_net_1 ), .B(
        \un1_next_int[4] ), .C(N333), .Y(N433));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I207_un1_Y_0 (.A(N508), .B(N539)
        , .Y(ADD_26x26_fast_I207_un1_Y_0));
    NOR3 inf_abs0_a_0_I_8 (.A(sr_new[0]), .B(sr_new[2]), .C(sr_new[1]), 
        .Y(N_11_0));
    AND3 inf_abs1_a_1_I_30 (.A(\DWACT_FINC_E_0[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E_0[6] ));
    MX2 \inf_abs1[3]  (.A(sr_old[3]), .B(\inf_abs1_a_1[3] ), .S(
        sr_old[12]), .Y(\inf_abs1[3]_net_1 ));
    XNOR2 inf_abs0_a_0_I_35 (.A(sr_new[12]), .B(N_2), .Y(
        \inf_abs0_a_0[12] ));
    NOR2 \state_RNIB3LN[1]  (.A(\state[0]_net_1 ), .B(\state[1]_net_1 )
        , .Y(N_46_1));
    OR2 \state_RNITN1H5[1]  (.A(\un18_next_int_m[10] ), .B(
        \inf_abs1_m[10] ), .Y(\un1_next_int_iv_0[10] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I188_Y (.A(N467), .B(I144_un1_Y), 
        .C(I188_un1_Y), .Y(N637));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I178_un1_Y (.A(N512), .B(N527), 
        .Y(I178_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I170_un1_Y (.A(N504), .B(N519), 
        .Y(I170_un1_Y));
    OR2 \state_RNIT6SR7[0]  (.A(\un1_next_int_iv_1[9] ), .B(
        \un2_next_int_m[9] ), .Y(\un1_next_int[9] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I45_Y (.A(integral[14]), .B(
        integral[15]), .C(\un1_next_int_0_iv_0[13] ), .Y(N413));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I137_Y (.A(N419), .B(N415), .C(
        N460), .Y(N514));
    XNOR2 inf_abs0_a_0_I_9 (.A(sr_new[3]), .B(N_11_0), .Y(
        \inf_abs0_a_0[3] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I3_P0N (.A(\un1_next_int_iv_0[3] )
        , .B(\un1_next_int_iv_1[3] ), .C(\integ[3]_net_1 ), .Y(N327));
    AX1D un1_integ_0_0_ADD_26x26_fast_I233_Y_0 (.A(
        \un1_next_int_iv_0[3] ), .B(\un1_next_int_iv_1[3] ), .C(
        \integ[3]_net_1 ), .Y(ADD_26x26_fast_I233_Y_0));
    NOR2B \state_RNO[0]  (.A(N_46_1), .B(calc_int), .Y(
        \state_RNO_7[0] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I50_Y (.A(I50_un1_Y), .B(N353), 
        .Y(N418));
    AO1 un1_integ_0_0_ADD_26x26_fast_I204_Y_3 (.A(N502), .B(N517), .C(
        ADD_26x26_fast_I204_Y_2), .Y(ADD_26x26_fast_I204_Y_3));
    XNOR2 inf_abs1_a_1_I_20 (.A(sr_old[7]), .B(N_7), .Y(
        \inf_abs1_a_1[7] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I74_un1_Y (.A(N318), .B(
        \un1_next_int[0] ), .Y(I74_un1_Y));
    OR2 \state_RNIS3I11_0[1]  (.A(next_int_1_sqmuxa), .B(
        next_int_0_sqmuxa_1), .Y(\un1_next_int_0_iv[13] ));
    OR3 \state_RNI5RGH8[0]  (.A(\inf_abs0_m[7] ), .B(
        \un1_next_int_iv_0[7] ), .C(\un2_next_int_m[7] ), .Y(
        \un1_next_int[7] ));
    OA1B un1_integ_0_0_ADD_26x26_fast_I36_Y (.A(integral[19]), .B(
        integral[18]), .C(\un1_next_int_0_iv_0[13] ), .Y(N404));
    NOR3A inf_abs1_a_1_I_31 (.A(\DWACT_FINC_E_0[6] ), .B(sr_old[9]), 
        .C(sr_old[10]), .Y(N_3_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I136_un1_Y (.A(N467), .B(N460), 
        .Y(I136_un1_Y));
    OR2 un1_integ_0_0_ADD_26x26_fast_I0_P0N (.A(N_3), .B(
        \integ[0]_net_1 ), .Y(N318));
    OR2 \state_RNIMLQF5[0]  (.A(\un1_next_int_iv_1[2] ), .B(
        \un1_next_int_iv_0[2] ), .Y(\un1_next_int[2] ));
    OR2 \state_RNIIMU77[0]  (.A(\un1_next_int_iv_1[6] ), .B(
        \inf_abs1_m[6] ), .Y(\un1_next_int[6] ));
    NOR2 inf_abs1_a_1_I_6 (.A(sr_old[0]), .B(sr_old[1]), .Y(N_12_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I55_Y (.A(N345), .B(N348), .Y(
        N423));
    OR2 \state_RNINO2D3[0]  (.A(\un1_next_int_iv_0[6] ), .B(
        \un2_next_int_m[6] ), .Y(\un1_next_int_iv_1[6] ));
    OA1 un1_integ_0_0_ADD_26x26_fast_I205_un1_Y (.A(N535), .B(
        I195_un1_Y), .C(ADD_26x26_fast_I205_un1_Y_0), .Y(I205_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I163_un1_Y (.A(N490), .B(
        \un1_next_int[0] ), .Y(I163_un1_Y));
    AO1 \state_RNI7F1S1[0]  (.A(sr_new[3]), .B(next_int_1_sqmuxa), .C(
        \un2_next_int_m[3] ), .Y(\un1_next_int_iv_1[3] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I120_un1_Y (.A(N439), .B(N442), 
        .Y(I120_un1_Y));
    NOR2 inf_abs1_a_1_I_21 (.A(sr_old[6]), .B(sr_old[7]), .Y(
        \DWACT_FINC_E[3] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I206_Y_1 (.A(N402), .B(N398), .C(
        N459), .Y(ADD_26x26_fast_I206_Y_1));
    OA1 un1_integ_0_0_ADD_26x26_fast_I5_G0N (.A(\un2_next_int_m[5] ), 
        .B(\un1_next_int_iv_1[5] ), .C(\integ[5]_net_1 ), .Y(N332));
    AND3 inf_abs0_a_0_I_24 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(
        \DWACT_FINC_E[4] ));
    DFN1E0C0 \integ[7]  (.D(\un1_integ[7] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(integral[7]));
    AO1 un1_integ_0_0_ADD_26x26_fast_I207_Y_2 (.A(
        ADD_26x26_fast_I207_un1_Y_0), .B(N524), .C(
        ADD_26x26_fast_I207_Y_1), .Y(ADD_26x26_fast_I207_Y_2));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I4_G0N (.A(\un1_next_int[4] ), 
        .B(\integ[4]_net_1 ), .Y(N329));
    OR2 un1_integ_0_0_ADD_26x26_fast_I195_Y (.A(N535), .B(I195_un1_Y), 
        .Y(N658));
    OA1 un1_integ_0_0_ADD_26x26_fast_I206_un1_Y_0 (.A(N483), .B(
        I160_un1_Y), .C(N506), .Y(ADD_26x26_fast_I206_un1_Y_0));
    NOR3B \state_RNIP0022[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0_a_0[12] ), .Y(\un2_next_int_m[12] ));
    XNOR2 inf_abs1_a_1_I_14 (.A(sr_old[5]), .B(N_9), .Y(
        \inf_abs1_a_1[5] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I234_Y (.A(N489), .B(I163_un1_Y), 
        .C(ADD_26x26_fast_I234_Y_0), .Y(\un1_integ[4] ));
    OR3 un1_integ_0_0_ADD_26x26_fast_I205_Y_2 (.A(N400), .B(
        ADD_26x26_fast_I205_Y_0), .C(N457), .Y(ADD_26x26_fast_I205_Y_2)
        );
    NOR2B un1_integ_0_0_ADD_26x26_fast_I174_un1_Y (.A(N508), .B(N523), 
        .Y(I174_un1_Y));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I162_un1_Y (.A(N488), .B(N442), 
        .Y(I162_un1_Y));
    AX1D un1_integ_0_0_ADD_26x26_fast_I240_Y (.A(N531), .B(I193_un1_Y), 
        .C(ADD_26x26_fast_I240_Y_0), .Y(\un1_integ[10] ));
    DFN1E0C0 \integ[8]  (.D(\un1_integ[8] ), .CLK(clk_c), .CLR(n_rst_c)
        , .E(N_46_1_0), .Q(integral[8]));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I85_Y (.A(N407), .B(N403), .Y(
        N456));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I251_Y_0 (.A(integral[21]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I251_Y_0));
    AO1 un1_integ_0_0_ADD_26x26_fast_I152_Y (.A(N483), .B(N476), .C(
        N475), .Y(N529));
    AND3 inf_abs0_a_0_I_22 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E_0[2] ), .C(\DWACT_FINC_E_0[3] ), .Y(N_6_0));
    OR2 un1_integ_0_0_ADD_26x26_fast_I9_P0N (.A(\un1_next_int[9] ), .B(
        integral[9]), .Y(N345));
    OA1 un1_integ_0_0_ADD_26x26_fast_I208_un1_Y_0 (.A(N487), .B(
        I162_un1_Y), .C(N510), .Y(ADD_26x26_fast_I208_un1_Y_0));
    NOR2B \state_RNIIHBH[0]  (.A(sr_new[8]), .B(next_int_1_sqmuxa), .Y(
        \inf_abs0_m[8] ));
    AO1B un1_integ_0_0_ADD_26x26_fast_I31_Y (.A(integral[22]), .B(
        integral[21]), .C(\un1_next_int_0_iv_0[13] ), .Y(N399));
    XNOR2 inf_abs1_a_1_I_12 (.A(sr_old[4]), .B(N_10_0), .Y(
        \inf_abs1_a_1[4] ));
    AX1D un1_integ_0_0_ADD_26x26_fast_I235_Y_0 (.A(\un2_next_int_m[5] )
        , .B(\un1_next_int_iv_1[5] ), .C(\integ[5]_net_1 ), .Y(
        ADD_26x26_fast_I235_Y_0));
    OR2 \state_RNIFGBI1[0]  (.A(\un18_next_int_m[4] ), .B(
        \inf_abs0_m[4] ), .Y(\un1_next_int_iv_0[4] ));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I56_un1_Y (.A(integral[8]), .B(
        \un1_next_int[8] ), .C(N345), .Y(I56_un1_Y));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I241_Y (.A(N649), .B(
        ADD_26x26_fast_I241_Y_0), .Y(\un1_integ[11] ));
    NOR3 inf_abs0_a_0_I_18 (.A(sr_new[4]), .B(sr_new[3]), .C(sr_new[5])
        , .Y(\DWACT_FINC_E_0[2] ));
    OR2 un1_integ_0_0_ADD_26x26_fast_I11_P0N (.A(\un1_next_int[11] ), 
        .B(integral[11]), .Y(N351));
    MX2 \inf_abs0[1]  (.A(sr_new[1]), .B(\inf_abs0_a_0[1] ), .S(
        sr_new_0_0), .Y(\inf_abs0[1]_net_1 ));
    XNOR2 un1_integ_0_0_ADD_26x26_fast_I243_Y_0 (.A(integral[13]), .B(
        \un1_next_int_0_iv[13] ), .Y(ADD_26x26_fast_I243_Y_0));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I105_Y (.A(N423), .B(N427), .Y(
        N476));
    MX2 \inf_abs0[11]  (.A(sr_new[11]), .B(\inf_abs0_a_0[11] ), .S(
        sr_new_0_0), .Y(\inf_abs0[11]_net_1 ));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I238_Y_0 (.A(\un1_next_int[8] ), 
        .B(integral[8]), .Y(ADD_26x26_fast_I238_Y_0));
    XOR2 inf_abs1_a_1_I_5 (.A(sr_old[0]), .B(sr_old[1]), .Y(
        \inf_abs1_a_1[1] ));
    NOR2B un1_integ_0_0_ADD_26x26_fast_I101_Y (.A(N419), .B(N423), .Y(
        N472));
    MAJ3 un1_integ_0_0_ADD_26x26_fast_I66_Y (.A(N326), .B(
        \integ[4]_net_1 ), .C(\un1_next_int[4] ), .Y(N434));
    AX1D un1_integ_0_0_ADD_26x26_fast_I248_Y (.A(
        ADD_26x26_fast_I211_Y_1), .B(ADD_26x26_fast_I211_Y_0), .C(
        ADD_26x26_fast_I248_Y_0), .Y(\un1_integ[18] ));
    AO1 \state_RNI3IGP3[1]  (.A(\inf_abs1[3]_net_1 ), .B(
        next_int_0_sqmuxa_1), .C(\un18_next_int_m[3] ), .Y(
        \un1_next_int_iv_0[3] ));
    NOR3B \state_RNI06J52[0]  (.A(sr_new[12]), .B(\state[0]_net_1 ), 
        .C(\inf_abs0[7]_net_1 ), .Y(\un2_next_int_m[7] ));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I99_Y (.A(N348), .B(N351), .C(
        N417), .Y(N470));
    OR2 un1_integ_0_0_ADD_26x26_fast_I92_Y (.A(N414), .B(N410), .Y(
        N463));
    OA1 un1_integ_0_0_ADD_26x26_fast_I191_un1_Y (.A(N489), .B(
        I163_un1_Y), .C(N528), .Y(I191_un1_Y));
    XA1A \state_RNIKB5M1[1]  (.A(sr_old[12]), .B(\inf_abs1[0]_net_1 ), 
        .C(\state[1]_net_1 ), .Y(\un1_next_int_iv_0[0] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I72_Y (.A(N317), .B(N321), .C(
        N320), .Y(N440));
    OA1B un1_integ_0_0_ADD_26x26_fast_I46_Y (.A(integral[13]), .B(
        integral[14]), .C(\un1_next_int_0_iv_0[13] ), .Y(N414));
    OR2 \state_RNI4PBS7[0]  (.A(\un1_next_int_iv_0[10] ), .B(
        \inf_abs0_m[10] ), .Y(\un1_next_int_iv_1[10] ));
    NOR3 inf_abs1_a_1_I_33 (.A(sr_old[10]), .B(sr_old[9]), .C(
        sr_old[11]), .Y(\DWACT_FINC_E_0[7] ));
    AO1 un1_integ_0_0_ADD_26x26_fast_I116_Y (.A(N438), .B(N435), .C(
        N434), .Y(N487));
    AO1 un1_integ_0_0_ADD_26x26_fast_I112_Y (.A(N434), .B(N431), .C(
        N430), .Y(N483));
    NOR2A inf_abs0_a_0_I_25 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .Y(
        N_5));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I213_un1_Y_0 (.A(N482), .B(N490)
        , .C(\un1_next_int[0] ), .Y(ADD_26x26_fast_I213_un1_Y_0));
    NOR3C un1_integ_0_0_ADD_26x26_fast_I210_un1_Y (.A(N530), .B(N491), 
        .C(N514), .Y(I210_un1_Y));
    XOR2 un1_integ_0_0_ADD_26x26_fast_I234_Y_0 (.A(\integ[4]_net_1 ), 
        .B(\un1_next_int[4] ), .Y(ADD_26x26_fast_I234_Y_0));
    NOR3A inf_abs0_a_0_I_27 (.A(\DWACT_FINC_E[4] ), .B(sr_new[8]), .C(
        sr_new[9]), .Y(N_4_0));
    
endmodule


module error_calc_13s_12s_4_3(
       cur_error,
       LED_15_i_0,
       LED_15,
       average,
       calc_error,
       n_rst_c,
       clk_c
    );
output [12:0] cur_error;
input  LED_15_i_0;
input  [7:0] LED_15;
input  [6:2] average;
input  calc_error;
input  n_rst_c;
input  clk_c;

    wire N_40, N_38, GND, VCC;
    
    AX1B un2_diffreg_1_m37 (.A(LED_15[5]), .B(LED_15[6]), .C(LED_15[7])
        , .Y(N_38));
    DFN1E1C0 \diffreg[3]  (.D(average[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[3]));
    XNOR2 un2_diffreg_1_m39 (.A(LED_15[6]), .B(LED_15[5]), .Y(N_40));
    VCC VCC_i (.Y(VCC));
    DFN1E1C0 \diffreg[7]  (.D(LED_15[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[7]));
    DFN1E1C0 \diffreg[1]  (.D(average[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[1]));
    DFN1E1C0 \diffreg[12]  (.D(N_38), .CLK(clk_c), .CLR(n_rst_c), .E(
        calc_error), .Q(cur_error[12]));
    DFN1E1C0 \diffreg[11]  (.D(N_40), .CLK(clk_c), .CLR(n_rst_c), .E(
        calc_error), .Q(cur_error[11]));
    GND GND_i (.Y(GND));
    DFN1E1C0 \diffreg[9]  (.D(LED_15[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[9]));
    DFN1E1C0 \diffreg[8]  (.D(LED_15[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[8]));
    DFN1E1C0 \diffreg[6]  (.D(LED_15[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[6]));
    DFN1E1C0 \diffreg[10]  (.D(LED_15_i_0), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[10]));
    DFN1E1C0 \diffreg[5]  (.D(LED_15[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[5]));
    DFN1E1C0 \diffreg[4]  (.D(average[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[4]));
    DFN1E1C0 \diffreg[2]  (.D(average[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[2]));
    DFN1E1C0 \diffreg[0]  (.D(average[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(calc_error), .Q(cur_error[0]));
    
endmodule


module derivative_calc_13s_4_3(
       derivative_0,
       sr_prev,
       sr_new,
       deriv_enable,
       n_rst_c,
       clk_c
    );
output derivative_0;
input  [12:0] sr_prev;
input  [12:0] sr_new;
input  deriv_enable;
input  n_rst_c;
input  clk_c;

    wire SUB_13x13_medium_area_I49_Y_1, N208, N176, 
        SUB_13x13_medium_area_I49_Y_0, 
        SUB_13x13_medium_area_I26_un1_Y_0, 
        SUB_13x13_medium_area_I49_un1_Y_1, 
        SUB_13x13_medium_area_I49_un1_Y_0, N_15, 
        SUB_13x13_medium_area_I42_Y_1, N218, N180, 
        SUB_13x13_medium_area_I42_Y_0, 
        SUB_13x13_medium_area_I30_un1_Y_0, 
        SUB_13x13_medium_area_I42_un1_Y_1, 
        SUB_13x13_medium_area_I42_un1_Y_0, N_7, 
        SUB_13x13_medium_area_I41_Y_0, 
        SUB_13x13_medium_area_I34_un1_Y_0, 
        SUB_13x13_medium_area_I41_un1_Y_0, N_5, 
        SUB_13x13_medium_area_I32_un1_Y_0, 
        SUB_13x13_medium_area_I28_un1_Y_0, N_24, N226, N204, N212, 
        N222, N185, N_21, N_13, GND, VCC;
    
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I34_un1_Y_0 (.A(
        sr_new[1]), .B(sr_prev[1]), .Y(
        SUB_13x13_medium_area_I34_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y_0 (.A(
        SUB_13x13_medium_area_I30_un1_Y_0), .B(sr_new[6]), .C(
        sr_prev[6]), .Y(SUB_13x13_medium_area_I42_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I15_S (.A(sr_prev[2]), 
        .B(sr_new[2]), .Y(N_5));
    OR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I36_Y (.A(sr_prev[0]), 
        .B(sr_new[0]), .Y(N185));
    XNOR3 un2_deriv_out_0_0_SUB_13x13_medium_area_I82_Y (.A(sr_new[12])
        , .B(sr_prev[12]), .C(N226), .Y(N_24));
    VCC VCC_i (.Y(VCC));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I64_Y (.A(N204), .B(
        sr_new[11]), .C(sr_prev[11]), .Y(N226));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I41_Y_0 (.A(
        SUB_13x13_medium_area_I34_un1_Y_0), .B(sr_new[2]), .C(
        sr_prev[2]), .Y(SUB_13x13_medium_area_I41_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I19_S (.A(sr_prev[6]), 
        .B(sr_new[6]), .Y(N_13));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I42_un1_Y_0 (.A(
        sr_new[4]), .B(sr_prev[4]), .C(N_7), .Y(
        SUB_13x13_medium_area_I42_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I28_Y (.A(
        SUB_13x13_medium_area_I28_un1_Y_0), .B(sr_new[8]), .C(
        sr_prev[8]), .Y(N208));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y_1 (.A(N218), .B(
        N180), .C(SUB_13x13_medium_area_I42_Y_0), .Y(
        SUB_13x13_medium_area_I42_Y_1));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I28_un1_Y_0 (.A(
        sr_new[7]), .B(sr_prev[7]), .Y(
        SUB_13x13_medium_area_I28_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y_0 (.A(
        SUB_13x13_medium_area_I26_un1_Y_0), .B(sr_new[10]), .C(
        sr_prev[10]), .Y(SUB_13x13_medium_area_I49_Y_0));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I20_S (.A(sr_prev[7]), 
        .B(sr_new[7]), .Y(N_15));
    DFN1E1C0 \deriv_out[12]  (.D(N_24), .CLK(clk_c), .CLR(n_rst_c), .E(
        deriv_enable), .Q(derivative_0));
    GND GND_i (.Y(GND));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I23_S (.A(sr_prev[10])
        , .B(sr_new[10]), .Y(N_21));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I26_un1_Y_0 (.A(
        sr_new[9]), .B(sr_prev[9]), .Y(
        SUB_13x13_medium_area_I26_un1_Y_0));
    AO13 un2_deriv_out_0_0_SUB_13x13_medium_area_I32_Y (.A(
        SUB_13x13_medium_area_I32_un1_Y_0), .B(sr_new[4]), .C(
        sr_prev[4]), .Y(N218));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I30_un1_Y_0 (.A(
        sr_new[5]), .B(sr_prev[5]), .Y(
        SUB_13x13_medium_area_I30_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y (.A(
        SUB_13x13_medium_area_I49_un1_Y_1), .B(N212), .C(
        SUB_13x13_medium_area_I49_Y_1), .Y(N204));
    NOR2A un2_deriv_out_0_0_SUB_13x13_medium_area_I32_un1_Y_0 (.A(
        sr_new[3]), .B(sr_prev[3]), .Y(
        SUB_13x13_medium_area_I32_un1_Y_0));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I31_Y (.A(sr_new[5]), 
        .B(sr_prev[5]), .C(N_13), .Y(N180));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I41_un1_Y_0 (.A(
        sr_new[1]), .B(sr_prev[1]), .C(N_5), .Y(
        SUB_13x13_medium_area_I41_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I49_Y_1 (.A(N208), .B(
        N176), .C(SUB_13x13_medium_area_I49_Y_0), .Y(
        SUB_13x13_medium_area_I49_Y_1));
    XOR2 un2_deriv_out_0_0_SUB_13x13_medium_area_I16_S (.A(sr_prev[3]), 
        .B(sr_new[3]), .Y(N_7));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I42_Y (.A(
        SUB_13x13_medium_area_I42_un1_Y_1), .B(N222), .C(
        SUB_13x13_medium_area_I42_Y_1), .Y(N212));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I27_Y (.A(sr_new[9]), 
        .B(sr_prev[9]), .C(N_21), .Y(N176));
    NOR2B un2_deriv_out_0_0_SUB_13x13_medium_area_I49_un1_Y_1 (.A(
        SUB_13x13_medium_area_I49_un1_Y_0), .B(N176), .Y(
        SUB_13x13_medium_area_I49_un1_Y_1));
    XA1C un2_deriv_out_0_0_SUB_13x13_medium_area_I49_un1_Y_0 (.A(
        sr_new[8]), .B(sr_prev[8]), .C(N_15), .Y(
        SUB_13x13_medium_area_I49_un1_Y_0));
    AO1 un2_deriv_out_0_0_SUB_13x13_medium_area_I41_Y (.A(
        SUB_13x13_medium_area_I41_un1_Y_0), .B(N185), .C(
        SUB_13x13_medium_area_I41_Y_0), .Y(N222));
    NOR2B un2_deriv_out_0_0_SUB_13x13_medium_area_I42_un1_Y_1 (.A(
        SUB_13x13_medium_area_I42_un1_Y_0), .B(N180), .Y(
        SUB_13x13_medium_area_I42_un1_Y_1));
    
endmodule


module pwm_tx_200s_32s_13s_10_1000000s_45s(
       off_div,
       act_ctl_5_0,
       pwm_chg,
       pwm_chg_0,
       n_rst_c,
       clk_c,
       act_ctl_5_8,
       act_ctl_5_7,
       act_ctl_5_2,
       act_ctl_5_4,
       act_ctl_5_3,
       primary_15_c
    );
input  [31:0] off_div;
input  act_ctl_5_0;
input  pwm_chg;
input  pwm_chg_0;
input  n_rst_c;
input  clk_c;
input  act_ctl_5_8;
input  act_ctl_5_7;
input  act_ctl_5_2;
input  act_ctl_5_4;
input  act_ctl_5_3;
output primary_15_c;

    wire N_403_0, I_140_8, I_140_7, \DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] , \DWACT_COMP0_E[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] , N_21, \counter[9]_net_1 , 
        N_7, \counter[3]_net_1 , N_10, N_17, N_13, \counter[8]_net_1 , 
        N_8, N_2, \counter[2]_net_1 , counter_63_0, 
        \counter[30]_net_1 , cur_pwm_RNI9RT933_0_net_1, 
        counter_m6_0_a2_7, counter_m6_0_a2_2, counter_m6_0_a2_1, 
        counter_m6_0_a2_6, \counter[16]_net_1 , \counter[18]_net_1 , 
        counter_m6_0_a2_4, \counter[15]_net_1 , \counter[10]_net_1 , 
        \counter[17]_net_1 , \counter[13]_net_1 , \counter[14]_net_1 , 
        \counter[11]_net_1 , \counter[12]_net_1 , counter_c18, 
        counter_c8, counter_n30, counter_c29, counter_n29, 
        \counter[29]_net_1 , counter_c28, counter_n28, counter_n28_tz, 
        \counter[27]_net_1 , counter_c26, \counter[28]_net_1 , 
        counter_n27, counter_n26, counter_n26_tz, \counter[25]_net_1 , 
        counter_c24, \counter[26]_net_1 , counter_n25, counter_n24, 
        counter_n24_tz, \counter[23]_net_1 , counter_c22, 
        \counter[24]_net_1 , counter_n23, counter_n22, counter_n22_tz, 
        \counter[21]_net_1 , counter_c20, \counter[22]_net_1 , 
        counter_n21, counter_n20, counter_n20_tz, \counter[19]_net_1 , 
        \counter[20]_net_1 , counter_n19, counter_n18, counter_c17, 
        counter_n17, counter_c16, counter_n16, counter_c15, 
        counter_n15, counter_c14, counter_n14, counter_c13, 
        counter_n13, counter_c12, counter_n12, counter_c11, 
        counter_n11, counter_c10, counter_n10, counter_n10_tz, 
        counter_n9, counter_n8, counter_n8_tz, \counter[7]_net_1 , 
        counter_c6, counter_n7, counter_n6, counter_n6_tz, 
        \counter[5]_net_1 , counter_c4, \counter[6]_net_1 , counter_n5, 
        counter_n4, counter_n4_tz, counter_c2, \counter[4]_net_1 , 
        counter_n3, counter_n2, counter_n2_tz, \counter[1]_net_1 , 
        \counter[0]_net_1 , \off_time[4] , \off_reg[4]_net_1 , 
        \off_time[9] , \off_reg[9]_net_1 , \off_time[10] , 
        \off_reg[10]_net_1 , \off_time[13] , \off_reg[13]_net_1 , 
        \off_time[14] , \off_reg[14]_net_1 , \off_time[19] , 
        \off_reg[19]_net_1 , \off_time[27] , \off_reg[27]_net_1 , 
        \off_time[15] , \off_reg[15]_net_1 , \off_time[22] , 
        \off_reg[22]_net_1 , \off_time[28] , \off_reg[28]_net_1 , 
        \off_time[16] , \off_reg[16]_net_1 , \off_time[11] , 
        \off_reg[11]_net_1 , \off_time[6] , \off_reg[6]_net_1 , 
        \off_time[24] , \off_reg[24]_net_1 , \off_time[29] , 
        \off_reg[29]_net_1 , \off_time[7] , \off_reg[7]_net_1 , 
        \off_time[17] , \off_reg[17]_net_1 , \off_time[18] , 
        \off_reg[18]_net_1 , \off_time[3] , \off_reg[3]_net_1 , 
        \off_time[23] , \off_reg[23]_net_1 , \off_time[20] , 
        \off_reg[20]_net_1 , \off_time[21] , \off_reg[21]_net_1 , 
        \off_time[26] , \off_reg[26]_net_1 , \off_time[25] , 
        \off_reg[25]_net_1 , \off_time[8] , \off_reg[8]_net_1 , 
        \off_time[2] , \off_reg[2]_net_1 , \off_time[1] , 
        \off_reg[1]_net_1 , \off_time[0] , \off_reg[0]_net_1 , 
        \off_time[31] , \off_reg[31]_net_1 , \off_time[5] , 
        \off_reg[5]_net_1 , \off_time[30] , \off_reg[30]_net_1 , 
        \off_time[12] , \off_reg[12]_net_1 , counter_n31, N_322, 
        counter_n1, \counter_RNO_3[0] , \counter[31]_net_1 , 
        cur_pwm_RNO_3, \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] , N_11, N_6, N_4, N_16, 
        N_18, N_12, N_14, \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] , \DWACT_BL_EQUAL_0_E[0] , 
        \DWACT_BL_EQUAL_0_E[1] , \DWACT_BL_EQUAL_0_E[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] , \DWACT_COMP0_E_0[1] , 
        \DWACT_COMP0_E_0[2] , \DWACT_COMP0_E[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] , N_11_0, N_10_0, N_9, 
        N_6_0, N_8_0, N_7_0, N_5, N_2_0, N_3, N_4_0, N_21_0, N_20, 
        N_19, N_16_0, N_18_0, N_17_0, N_15, N_12_0, N_13_0, N_14_0, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] , 
        \DWACT_BL_EQUAL_0_E[4] , \DWACT_BL_EQUAL_0_E[3] , 
        \DWACT_BL_EQUAL_0_E_0[0] , \DWACT_BL_EQUAL_0_E_0[1] , 
        \DWACT_BL_EQUAL_0_E_0[2] , \DWACT_CMPLE_PO0_DWACT_COMP0_E[1] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[0] , N_31, N_30, N_29, N_26, 
        N_28, N_27, N_25, N_22, N_23, N_24, \ACT_LT4_E[3] , 
        \ACT_LT4_E[6] , \ACT_LT4_E[10] , \ACT_LT4_E[7] , 
        \ACT_LT4_E[8] , \ACT_LT4_E[5] , \ACT_LT4_E[4] , \ACT_LT4_E[0] , 
        \ACT_LT4_E[1] , \ACT_LT4_E[2] , \DWACT_BL_EQUAL_0_E_0[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] , 
        \DWACT_BL_EQUAL_0_E_1[0] , \DWACT_BL_EQUAL_0_E_1[1] , 
        \DWACT_BL_EQUAL_0_E_1[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] , 
        \DWACT_BL_EQUAL_0_E_2[0] , \DWACT_BL_EQUAL_0_E_2[1] , 
        \DWACT_BL_EQUAL_0_E_2[2] , \DWACT_BL_EQUAL_0_E_1[3] , 
        \DWACT_BL_EQUAL_0_E_0[4] , \DWACT_BL_EQUAL_0_E[5] , 
        \DWACT_BL_EQUAL_0_E[6] , \DWACT_BL_EQUAL_0_E[7] , 
        \DWACT_BL_EQUAL_0_E[8] , \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] , N_41, N_40, N_39, N_36, 
        N_38, N_37, N_35, N_32, N_33, N_34, \ACT_LT3_E[3] , 
        \ACT_LT3_E[4] , \ACT_LT3_E[5] , \ACT_LT3_E[0] , \ACT_LT3_E[1] , 
        \ACT_LT3_E[2] , \DWACT_BL_EQUAL_0_E_3[2] , 
        \DWACT_BL_EQUAL_0_E_3[1] , \DWACT_BL_EQUAL_0_E_3[0] , N_51, 
        N_50, N_49, N_46, N_48, N_47, N_45, N_42, N_43, N_44, 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] , 
        \DWACT_BL_EQUAL_0_E_1[4] , \DWACT_BL_EQUAL_0_E_2[3] , 
        \DWACT_BL_EQUAL_0_E_4[0] , \DWACT_BL_EQUAL_0_E_4[1] , 
        \DWACT_BL_EQUAL_0_E_4[2] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] , 
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] , 
        \DWACT_BL_EQUAL_0_E[12] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] , 
        \DWACT_BL_EQUAL_0_E_5[0] , \DWACT_BL_EQUAL_0_E_5[1] , 
        \DWACT_BL_EQUAL_0_E_5[2] , \DWACT_BL_EQUAL_0_E_3[3] , 
        \DWACT_BL_EQUAL_0_E_2[4] , \DWACT_BL_EQUAL_0_E_0[5] , 
        \DWACT_BL_EQUAL_0_E_0[6] , \DWACT_BL_EQUAL_0_E_0[7] , 
        \DWACT_BL_EQUAL_0_E_0[8] , \DWACT_BL_EQUAL_0_E[9] , 
        \DWACT_BL_EQUAL_0_E[10] , \DWACT_BL_EQUAL_0_E[11] , GND, VCC;
    
    DFN1C0 \counter[19]  (.D(counter_n19), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[19]_net_1 ));
    AND3 un1_counter_0_I_78 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] ));
    NOR3 un1_counter_2_0_I_17 (.A(\counter[20]_net_1 ), .B(
        \counter[19]_net_1 ), .C(\counter[21]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] ));
    AND2A un1_counter_0_I_51 (.A(\off_time[26] ), .B(
        \counter[26]_net_1 ), .Y(\ACT_LT3_E[5] ));
    NOR2A \off_reg_RNIRJ0K[24]  (.A(\off_reg[24]_net_1 ), .B(
        act_ctl_5_8), .Y(\off_time[24] ));
    DFN1E1C0 \off_reg[28]  (.D(off_div[28]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[28]_net_1 ));
    AX1C \counter_RNO_0[2]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .C(\counter[2]_net_1 ), .Y(counter_n2_tz));
    DFN1C0 \counter[28]  (.D(counter_n28), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[28]_net_1 ));
    XNOR2 un1_counter_0_I_73 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .Y(\DWACT_BL_EQUAL_0_E_2[2] ));
    OA1A un1_counter_0_I_136 (.A(N_6_0), .B(N_8_0), .C(N_7_0), .Y(
        N_11_0));
    OR2 un1_counter_2_0_I_116 (.A(\counter[6]_net_1 ), .B(act_ctl_5_3), 
        .Y(N_12));
    OA1A un1_counter_0_I_132 (.A(\counter[3]_net_1 ), .B(\off_time[3] )
        , .C(N_3), .Y(N_7_0));
    DFN1E1C0 \off_reg[15]  (.D(off_div[15]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[15]_net_1 ));
    DFN1E1C0 \off_reg[26]  (.D(off_div[26]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[26]_net_1 ));
    AND3 un1_counter_0_I_14 (.A(\DWACT_BL_EQUAL_0_E[9] ), .B(
        \DWACT_BL_EQUAL_0_E[10] ), .C(\DWACT_BL_EQUAL_0_E[11] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] ));
    XA1B \counter_RNO[11]  (.A(\counter[11]_net_1 ), .B(counter_c10), 
        .C(N_403_0), .Y(counter_n11));
    DFN1C0 \counter[29]  (.D(counter_n29), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[29]_net_1 ));
    DFN1E1C0 \off_reg[5]  (.D(off_div[5]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[5]_net_1 ));
    NOR3 un1_counter_2_0_I_77 (.A(\counter[12]_net_1 ), .B(
        \counter[10]_net_1 ), .C(\counter[11]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] ));
    XNOR2 un1_counter_0_I_82 (.A(\counter[15]_net_1 ), .B(
        \off_time[15] ), .Y(\DWACT_BL_EQUAL_0_E_1[0] ));
    DFN1C0 \counter[11]  (.D(counter_n11), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[11]_net_1 ));
    XNOR2 un1_counter_0_I_109 (.A(\counter[6]_net_1 ), .B(
        \off_time[6] ), .Y(\DWACT_BL_EQUAL_0_E_0[1] ));
    OR2 \off_reg_RNISHSI[17]  (.A(\off_reg[17]_net_1 ), .B(act_ctl_5_7)
        , .Y(\off_time[17] ));
    NOR2B \counter_RNIF23M[11]  (.A(\counter[11]_net_1 ), .B(
        \counter[12]_net_1 ), .Y(counter_m6_0_a2_1));
    NOR2A un1_counter_2_0_I_118 (.A(act_ctl_5_3), .B(
        \counter[5]_net_1 ), .Y(N_14));
    OR2A un1_counter_0_I_103 (.A(\counter[14]_net_1 ), .B(
        \off_time[14] ), .Y(N_29));
    NOR2A \off_reg_RNIOH1K[30]  (.A(\off_reg[30]_net_1 ), .B(
        act_ctl_5_8), .Y(\off_time[30] ));
    NOR2A \counter_RNO[28]  (.A(counter_n28_tz), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n28));
    XA1B \counter_RNO[15]  (.A(\counter[15]_net_1 ), .B(counter_c14), 
        .C(N_403_0), .Y(counter_n15));
    XNOR2 un1_counter_0_I_25 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .Y(\DWACT_BL_EQUAL_0_E_2[3] ));
    NOR2B \counter_RNIJ63M[13]  (.A(\counter[13]_net_1 ), .B(
        \counter[14]_net_1 ), .Y(counter_m6_0_a2_2));
    AND2 un1_counter_0_I_114 (.A(\DWACT_BL_EQUAL_0_E[4] ), .B(
        \DWACT_BL_EQUAL_0_E[3] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] ));
    XNOR2 un1_counter_0_I_11 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .Y(\DWACT_BL_EQUAL_0_E_3[3] ));
    NOR2A \off_reg_RNIUM0K[27]  (.A(\off_reg[27]_net_1 ), .B(
        act_ctl_5_8), .Y(\off_time[27] ));
    AX1C \counter_RNO_0[22]  (.A(\counter[21]_net_1 ), .B(counter_c20), 
        .C(\counter[22]_net_1 ), .Y(counter_n22_tz));
    XA1B \counter_RNO[7]  (.A(\counter[7]_net_1 ), .B(counter_c6), .C(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n7));
    OA1A un1_counter_2_0_I_125 (.A(N_16), .B(N_18), .C(N_17), .Y(N_21));
    DFN1E1C0 \off_reg[2]  (.D(off_div[2]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[2]_net_1 ));
    XNOR2 un1_counter_0_I_72 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .Y(\DWACT_BL_EQUAL_0_E_1[3] ));
    OA1 un1_counter_0_I_126 (.A(N_21_0), .B(N_20), .C(N_19), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] ));
    DFN1C0 \counter[6]  (.D(counter_n6), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[6]_net_1 ));
    AO1C un1_counter_0_I_122 (.A(\counter[7]_net_1 ), .B(\off_time[7] )
        , .C(N_12_0), .Y(N_18_0));
    AX1C \counter_RNO[31]  (.A(counter_c29), .B(counter_63_0), .C(
        N_322), .Y(counter_n31));
    NOR3C \counter_RNIR7IOA[27]  (.A(\counter[27]_net_1 ), .B(
        counter_c26), .C(\counter[28]_net_1 ), .Y(counter_c28));
    DFN1C0 \counter[21]  (.D(counter_n21), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[21]_net_1 ));
    AND2 un1_counter_0_I_20 (.A(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] ), .B(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] ), .Y(
        \DWACT_COMP0_E_0[1] ));
    XOR2 un1_counter_2_0_I_109 (.A(act_ctl_5_3), .B(\counter[6]_net_1 )
        , .Y(\DWACT_BL_EQUAL_0_E[1] ));
    DFN1C0 \counter[3]  (.D(counter_n3), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[3]_net_1 ));
    DFN1C0 \counter[2]  (.D(counter_n2), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[2]_net_1 ));
    AND3 un1_counter_0_I_45 (.A(\DWACT_BL_EQUAL_0_E_3[2] ), .B(
        \DWACT_BL_EQUAL_0_E_3[1] ), .C(\DWACT_BL_EQUAL_0_E_3[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] ));
    NOR2A \off_reg_RNI4D43[5]  (.A(\off_reg[5]_net_1 ), .B(act_ctl_5_2)
        , .Y(\off_time[5] ));
    DFN1E1C0 \off_reg[23]  (.D(off_div[23]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[23]_net_1 ));
    NOR2A \counter_RNO[8]  (.A(counter_n8_tz), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n8));
    NOR2A un1_counter_2_0_I_121 (.A(N_13), .B(\counter[8]_net_1 ), .Y(
        N_17));
    XA1B \counter_RNO[13]  (.A(\counter[13]_net_1 ), .B(counter_c12), 
        .C(N_403_0), .Y(counter_n13));
    AO1C un1_counter_0_I_57 (.A(\off_time[20] ), .B(
        \counter[20]_net_1 ), .C(N_34), .Y(N_36));
    NOR3C \counter_RNIGR1M8[22]  (.A(\counter[21]_net_1 ), .B(
        counter_c20), .C(\counter[22]_net_1 ), .Y(counter_c22));
    DFN1E1C0 \off_reg[9]  (.D(off_div[9]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[9]_net_1 ));
    XNOR2 un1_counter_0_I_26 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(\DWACT_BL_EQUAL_0_E_4[2] ));
    AX1C \counter_RNO_0[4]  (.A(\counter[3]_net_1 ), .B(counter_c2), 
        .C(\counter[4]_net_1 ), .Y(counter_n4_tz));
    AO1C un1_counter_0_I_35 (.A(\off_time[28] ), .B(
        \counter[28]_net_1 ), .C(N_44), .Y(N_46));
    AO1 un1_counter_0_I_65 (.A(\DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] ), 
        .B(\DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] ), .C(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] ), .Y(\DWACT_COMP0_E[0] ));
    NOR2A un1_counter_2_0_I_135 (.A(act_ctl_5_4), .B(
        \counter[3]_net_1 ), .Y(N_10));
    NOR2B \counter_RNIERKJ6[16]  (.A(counter_c15), .B(
        \counter[16]_net_1 ), .Y(counter_c16));
    AND2 un1_counter_0_I_84 (.A(\DWACT_BL_EQUAL_0_E_0[3] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[1] ));
    NOR2A \off_reg_RNIODSI[13]  (.A(\off_reg[13]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[13] ));
    DFN1C0 cur_pwm (.D(cur_pwm_RNO_3), .CLK(clk_c), .CLR(n_rst_c), .Q(
        primary_15_c));
    XA1B \counter_RNO[12]  (.A(\counter[12]_net_1 ), .B(counter_c11), 
        .C(N_403_0), .Y(counter_n12));
    AOI1A un1_counter_0_I_95 (.A(\ACT_LT4_E[3] ), .B(\ACT_LT4_E[6] ), 
        .C(\ACT_LT4_E[10] ), .Y(\DWACT_CMPLE_PO0_DWACT_COMP0_E[0] ));
    OA1A un1_counter_0_I_40 (.A(N_46), .B(N_48), .C(N_47), .Y(N_51));
    XA1B \counter_RNO[1]  (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(N_403_0), .Y(counter_n1));
    NOR2B \counter_RNITSFI5[13]  (.A(counter_c12), .B(
        \counter[13]_net_1 ), .Y(counter_c13));
    DFN1C0 \counter[17]  (.D(counter_n17), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[17]_net_1 ));
    NOR2 un1_counter_2_0_I_129 (.A(\counter[0]_net_1 ), .B(act_ctl_5_3)
        , .Y(N_4));
    DFN1C0 \counter[4]  (.D(counter_n4), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[4]_net_1 ));
    AO1B un1_counter_2_0_I_131 (.A(act_ctl_5_0), .B(\counter[1]_net_1 )
        , .C(N_4), .Y(N_6));
    AND2 un1_counter_0_I_30 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[1] ));
    OR2A un1_counter_0_I_60 (.A(\counter[23]_net_1 ), .B(
        \off_time[23] ), .Y(N_39));
    DFN1E1C0 \off_reg[11]  (.D(off_div[11]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[11]_net_1 ));
    AND2 un1_counter_0_I_29 (.A(\DWACT_BL_EQUAL_0_E_1[4] ), .B(
        \DWACT_BL_EQUAL_0_E_2[3] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[1] ));
    DFN1E1C0 \off_reg[22]  (.D(off_div[22]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[22]_net_1 ));
    DFN1C0 \counter[10]  (.D(counter_n10), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[10]_net_1 ));
    NOR2A un1_counter_2_0_I_19 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] ), .B(\counter[31]_net_1 )
        , .Y(\DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] ));
    NOR2A un1_counter_0_I_46 (.A(\off_time[24] ), .B(
        \counter[24]_net_1 ), .Y(\ACT_LT3_E[0] ));
    GND GND_i (.Y(GND));
    DFN1C0 \counter[13]  (.D(counter_n13), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[13]_net_1 ));
    XNOR2 un1_counter_0_I_81 (.A(\counter[16]_net_1 ), .B(
        \off_time[16] ), .Y(\DWACT_BL_EQUAL_0_E_1[1] ));
    NOR2A un1_counter_0_I_90 (.A(\off_time[18] ), .B(
        \counter[18]_net_1 ), .Y(\ACT_LT4_E[5] ));
    XNOR2 un1_counter_0_I_74 (.A(\counter[11]_net_1 ), .B(
        \off_time[11] ), .Y(\DWACT_BL_EQUAL_0_E_2[1] ));
    NOR2B un1_counter_2_0_I_140 (.A(\DWACT_COMP0_E[2] ), .B(
        \DWACT_COMP0_E[1] ), .Y(I_140_7));
    OA1A un1_counter_0_I_36 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .C(N_43), .Y(N_47));
    XNOR2 un1_counter_0_I_66 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\DWACT_BL_EQUAL_0_E[8] ));
    AND3 un1_counter_0_I_17 (.A(\DWACT_BL_EQUAL_0_E_5[0] ), .B(
        \DWACT_BL_EQUAL_0_E_5[1] ), .C(\DWACT_BL_EQUAL_0_E_5[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] ));
    DFN1E1C0 \off_reg[17]  (.D(off_div[17]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[17]_net_1 ));
    NOR3C \counter_RNI9AO97[9]  (.A(\counter[9]_net_1 ), .B(counter_c8)
        , .C(counter_m6_0_a2_7), .Y(counter_c18));
    AX1C \counter_RNO_0[10]  (.A(\counter[9]_net_1 ), .B(counter_c8), 
        .C(\counter[10]_net_1 ), .Y(counter_n10_tz));
    DFN1C0 \counter[12]  (.D(counter_n12), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[12]_net_1 ));
    OR2A un1_counter_0_I_130 (.A(\off_time[4] ), .B(\counter[4]_net_1 )
        , .Y(N_5));
    NOR2B un1_counter_2_0_I_139 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E[2] )
        , .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ), .Y(
        \DWACT_COMP0_E[2] ));
    NOR2A \off_reg_RNI7G43[8]  (.A(\off_reg[8]_net_1 ), .B(act_ctl_5_2)
        , .Y(\off_time[8] ));
    DFN1C0 \counter[27]  (.D(counter_n27), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[27]_net_1 ));
    OR2A un1_counter_0_I_96 (.A(\off_time[11] ), .B(
        \counter[11]_net_1 ), .Y(N_22));
    NOR3C \counter_RNIO20U2[5]  (.A(\counter[5]_net_1 ), .B(counter_c4)
        , .C(\counter[6]_net_1 ), .Y(counter_c6));
    AOI1A un1_counter_0_I_49 (.A(\ACT_LT3_E[0] ), .B(\ACT_LT3_E[1] ), 
        .C(\ACT_LT3_E[2] ), .Y(\ACT_LT3_E[3] ));
    NOR2B \counter_RNINGHT5[14]  (.A(counter_c13), .B(
        \counter[14]_net_1 ), .Y(counter_c14));
    AX1C \counter_RNO_0[20]  (.A(\counter[19]_net_1 ), .B(counter_c18), 
        .C(\counter[20]_net_1 ), .Y(counter_n20_tz));
    DFN1C0 \counter[20]  (.D(counter_n20), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[20]_net_1 ));
    OA1A un1_counter_0_I_101 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .C(N_23), .Y(N_27));
    DFN1E1C0 \off_reg[19]  (.D(off_div[19]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[19]_net_1 ));
    XNOR2 un1_counter_0_I_71 (.A(\counter[10]_net_1 ), .B(
        \off_time[10] ), .Y(\DWACT_BL_EQUAL_0_E_2[0] ));
    OR2A un1_counter_0_I_116 (.A(\off_time[6] ), .B(\counter[6]_net_1 )
        , .Y(N_12_0));
    AO1C un1_counter_0_I_39 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .C(N_45), .Y(N_50));
    XA1B \counter_RNO[17]  (.A(\counter[17]_net_1 ), .B(counter_c16), 
        .C(N_403_0), .Y(counter_n17));
    XNOR2 un1_counter_0_I_69 (.A(\counter[16]_net_1 ), .B(
        \off_time[16] ), .Y(\DWACT_BL_EQUAL_0_E[6] ));
    XNOR2 un1_counter_0_I_112 (.A(\counter[9]_net_1 ), .B(
        \off_time[9] ), .Y(\DWACT_BL_EQUAL_0_E[4] ));
    OA1A un1_counter_0_I_105 (.A(N_26), .B(N_28), .C(N_27), .Y(N_31));
    DFN1C0 \counter[23]  (.D(counter_n23), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[23]_net_1 ));
    XA1B \counter_RNO[29]  (.A(\counter[29]_net_1 ), .B(counter_c28), 
        .C(N_403_0), .Y(counter_n29));
    NOR2A \off_reg_RNIMCTI[20]  (.A(\off_reg[20]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[20] ));
    NOR2A \off_reg_RNI6F43[7]  (.A(\off_reg[7]_net_1 ), .B(act_ctl_5_2)
        , .Y(\off_time[7] ));
    DFN1E1C0 \off_reg[25]  (.D(off_div[25]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[25]_net_1 ));
    NOR2B \counter_RNO_0[18]  (.A(counter_c16), .B(\counter[17]_net_1 )
        , .Y(counter_c17));
    DFN1C0 \counter[22]  (.D(counter_n22), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[22]_net_1 ));
    DFN1C0 \counter[15]  (.D(counter_n15), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[15]_net_1 ));
    AO1 un1_counter_0_I_107 (.A(\DWACT_CMPLE_PO0_DWACT_COMP0_E[1] ), 
        .B(\DWACT_CMPLE_PO0_DWACT_COMP0_E[2] ), .C(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] ));
    OR2A un1_counter_0_I_99 (.A(\off_time[14] ), .B(
        \counter[14]_net_1 ), .Y(N_25));
    OAI1 un1_counter_2_0_I_122 (.A(act_ctl_5_0), .B(\counter[7]_net_1 )
        , .C(N_12), .Y(N_18));
    AND2 un1_counter_2_0_I_115 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] ));
    OR2 \off_reg_RNIPESI[14]  (.A(\off_reg[14]_net_1 ), .B(act_ctl_5_7)
        , .Y(\off_time[14] ));
    XNOR2 un1_counter_0_I_108 (.A(\counter[5]_net_1 ), .B(
        \off_time[5] ), .Y(\DWACT_BL_EQUAL_0_E_0[0] ));
    NOR3C \counter_RNI3F432[4]  (.A(\counter[3]_net_1 ), .B(counter_c2)
        , .C(\counter[4]_net_1 ), .Y(counter_c4));
    NOR2A \off_reg_RNI0P0K[29]  (.A(\off_reg[29]_net_1 ), .B(
        act_ctl_5_8), .Y(\off_time[29] ));
    AX1C \counter_RNO_0[8]  (.A(\counter[7]_net_1 ), .B(counter_c6), 
        .C(\counter[8]_net_1 ), .Y(counter_n8_tz));
    AX1C \counter_RNO_0[28]  (.A(\counter[27]_net_1 ), .B(counter_c26), 
        .C(\counter[28]_net_1 ), .Y(counter_n28_tz));
    VCC VCC_i (.Y(VCC));
    AO1C un1_counter_0_I_120 (.A(\off_time[6] ), .B(\counter[6]_net_1 )
        , .C(N_14_0), .Y(N_16_0));
    DFN1E1C0 \off_reg[31]  (.D(off_div[31]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[31]_net_1 ));
    XA1B \counter_RNO[14]  (.A(\counter[14]_net_1 ), .B(counter_c13), 
        .C(N_403_0), .Y(counter_n14));
    XOR2 un1_counter_2_0_I_111 (.A(act_ctl_5_3), .B(\counter[7]_net_1 )
        , .Y(\DWACT_BL_EQUAL_0_E[2] ));
    DFN1E1C0 \off_reg[7]  (.D(off_div[7]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[7]_net_1 ));
    DFN1C0 \counter[1]  (.D(counter_n1), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[1]_net_1 ));
    XNOR2 un1_counter_0_I_2 (.A(\counter[19]_net_1 ), .B(
        \off_time[19] ), .Y(\DWACT_BL_EQUAL_0_E_5[0] ));
    NOR2A \counter_RNO[26]  (.A(counter_n26_tz), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n26));
    NOR2A un1_counter_0_I_55 (.A(\off_time[19] ), .B(
        \counter[19]_net_1 ), .Y(N_34));
    AO1 un1_counter_0_I_139 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_1[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_0[0] ), .Y(\DWACT_COMP0_E_0[2] )
        );
    XA1B \counter_RNO[5]  (.A(\counter[5]_net_1 ), .B(counter_c4), .C(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n5));
    AO1C un1_counter_0_I_133 (.A(\counter[2]_net_1 ), .B(\off_time[2] )
        , .C(N_2_0), .Y(N_8_0));
    OR2A un1_counter_2_0_I_132 (.A(\counter[3]_net_1 ), .B(act_ctl_5_3)
        , .Y(N_7));
    MX2C cur_pwm_RNI9RT933_0 (.A(I_140_8), .B(I_140_7), .S(
        primary_15_c), .Y(cur_pwm_RNI9RT933_0_net_1));
    DFN1C0 \counter[25]  (.D(counter_n25), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[25]_net_1 ));
    AND2A un1_counter_0_I_87 (.A(\off_time[16] ), .B(
        \counter[16]_net_1 ), .Y(\ACT_LT4_E[2] ));
    XA1B \counter_RNO[3]  (.A(\counter[3]_net_1 ), .B(counter_c2), .C(
        N_403_0), .Y(counter_n3));
    DFN1E1C0 \off_reg[6]  (.D(off_div[6]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[6]_net_1 ));
    AND3 un1_counter_0_I_28 (.A(\DWACT_BL_EQUAL_0_E_4[0] ), .B(
        \DWACT_BL_EQUAL_0_E_4[1] ), .C(\DWACT_BL_EQUAL_0_E_4[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[0] ));
    OR2A un1_counter_0_I_50 (.A(\off_time[26] ), .B(
        \counter[26]_net_1 ), .Y(\ACT_LT3_E[4] ));
    DFN1C0 \counter[5]  (.D(counter_n5), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[5]_net_1 ));
    MX2A cur_pwm_RNO (.A(I_140_8), .B(I_140_7), .S(primary_15_c), .Y(
        cur_pwm_RNO_3));
    XNOR2 un1_counter_0_I_4 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(\DWACT_BL_EQUAL_0_E[10] ));
    XNOR2 un1_counter_0_I_23 (.A(\counter[27]_net_1 ), .B(
        \off_time[27] ), .Y(\DWACT_BL_EQUAL_0_E_4[0] ));
    NOR3C \counter_RNI898N1[18]  (.A(\counter[16]_net_1 ), .B(
        \counter[18]_net_1 ), .C(counter_m6_0_a2_4), .Y(
        counter_m6_0_a2_6));
    NOR2A \counter_RNO[10]  (.A(counter_n10_tz), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n10));
    AND3 un1_counter_0_I_77 (.A(\DWACT_BL_EQUAL_0_E_2[0] ), .B(
        \DWACT_BL_EQUAL_0_E_2[1] ), .C(\DWACT_BL_EQUAL_0_E_2[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_4[0] ));
    XNOR2 un1_counter_0_I_3 (.A(\counter[30]_net_1 ), .B(
        \off_time[30] ), .Y(\DWACT_BL_EQUAL_0_E[11] ));
    XA1B \counter_RNO[21]  (.A(\counter[21]_net_1 ), .B(counter_c20), 
        .C(N_403_0), .Y(counter_n21));
    XNOR2 un1_counter_0_I_6 (.A(\counter[20]_net_1 ), .B(
        \off_time[20] ), .Y(\DWACT_BL_EQUAL_0_E_5[1] ));
    OR2A un1_counter_0_I_56 (.A(\off_time[23] ), .B(
        \counter[23]_net_1 ), .Y(N_35));
    AX1C \counter_RNO_0[24]  (.A(\counter[23]_net_1 ), .B(counter_c22), 
        .C(\counter[24]_net_1 ), .Y(counter_n24_tz));
    AND3 un1_counter_0_I_15 (.A(\DWACT_BL_EQUAL_0_E_0[6] ), .B(
        \DWACT_BL_EQUAL_0_E_0[7] ), .C(\DWACT_BL_EQUAL_0_E_0[8] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] ));
    AND2A un1_counter_0_I_48 (.A(\off_time[25] ), .B(
        \counter[25]_net_1 ), .Y(\ACT_LT3_E[2] ));
    NOR2A un1_counter_0_I_129 (.A(\off_time[0] ), .B(
        \counter[0]_net_1 ), .Y(N_4_0));
    XNOR2 un1_counter_0_I_9 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(\DWACT_BL_EQUAL_0_E[12] ));
    AO1 un1_counter_0_I_140 (.A(\DWACT_COMP0_E_0[1] ), .B(
        \DWACT_COMP0_E_0[2] ), .C(\DWACT_COMP0_E[0] ), .Y(I_140_8));
    OR2A un1_counter_0_I_123 (.A(\counter[9]_net_1 ), .B(\off_time[9] )
        , .Y(N_19));
    DFN1C0 \counter[16]  (.D(counter_n16), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[16]_net_1 ));
    OR2A un1_counter_0_I_38 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(N_49));
    XA1B \counter_RNO[25]  (.A(\counter[25]_net_1 ), .B(counter_c24), 
        .C(N_403_0), .Y(counter_n25));
    XNOR2 un1_counter_0_I_68 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\DWACT_BL_EQUAL_0_E[7] ));
    NOR2A \counter_RNO_0[31]  (.A(\counter[30]_net_1 ), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_63_0));
    NOR3C \counter_RNIER411[10]  (.A(\counter[15]_net_1 ), .B(
        \counter[10]_net_1 ), .C(\counter[17]_net_1 ), .Y(
        counter_m6_0_a2_4));
    XNOR2 un1_counter_0_I_43 (.A(\counter[25]_net_1 ), .B(
        \off_time[25] ), .Y(\DWACT_BL_EQUAL_0_E_3[1] ));
    AO1C un1_counter_0_I_59 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .C(N_32), .Y(N_38));
    DFN1E1C0 \off_reg[21]  (.D(off_div[21]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[21]_net_1 ));
    AO1C un1_counter_0_I_104 (.A(\counter[13]_net_1 ), .B(
        \off_time[13] ), .C(N_25), .Y(N_30));
    NOR2A \off_reg_RNILASI[10]  (.A(\off_reg[10]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[10] ));
    OR2 un1_counter_2_0_I_127 (.A(\counter[1]_net_1 ), .B(act_ctl_5_3), 
        .Y(N_2));
    XNOR2 un1_counter_0_I_10 (.A(\counter[24]_net_1 ), .B(
        \off_time[24] ), .Y(\DWACT_BL_EQUAL_0_E_0[5] ));
    NOR2A un1_counter_0_I_98 (.A(\off_time[10] ), .B(
        \counter[10]_net_1 ), .Y(N_24));
    NOR2A un1_counter_0_I_33 (.A(\off_time[27] ), .B(
        \counter[27]_net_1 ), .Y(N_44));
    OA1 un1_counter_0_I_63 (.A(N_41), .B(N_40), .C(N_39), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] ));
    NOR2A \off_reg_RNITL0K[26]  (.A(\off_reg[26]_net_1 ), .B(
        act_ctl_5_8), .Y(\off_time[26] ));
    NOR2A \counter_RNO[6]  (.A(counter_n6_tz), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n6));
    XA1B \counter_RNO[30]  (.A(\counter[30]_net_1 ), .B(counter_c29), 
        .C(N_403_0), .Y(counter_n30));
    XNOR2 un1_counter_0_I_110 (.A(\counter[8]_net_1 ), .B(
        \off_time[8] ), .Y(\DWACT_BL_EQUAL_0_E[3] ));
    DFN1E1C0 \off_reg[27]  (.D(off_div[27]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[27]_net_1 ));
    AND3 un1_counter_0_I_16 (.A(\DWACT_BL_EQUAL_0_E_3[3] ), .B(
        \DWACT_BL_EQUAL_0_E_2[4] ), .C(\DWACT_BL_EQUAL_0_E_0[5] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] ));
    OR2A un1_counter_0_I_93 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\ACT_LT4_E[8] ));
    DFN1E1C0 \off_reg[8]  (.D(off_div[8]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[8]_net_1 ));
    NOR3C \counter_RNIIV881[2]  (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .C(\counter[2]_net_1 ), .Y(counter_c2));
    DFN1C0 \counter[26]  (.D(counter_n26), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[26]_net_1 ));
    OR2 \off_reg_RNIRGSI[16]  (.A(\off_reg[16]_net_1 ), .B(act_ctl_5_7)
        , .Y(\off_time[16] ));
    XA1B \counter_RNO[23]  (.A(\counter[23]_net_1 ), .B(counter_c22), 
        .C(N_403_0), .Y(counter_n23));
    OA1B un1_counter_2_0_I_137 (.A(N_10), .B(N_11), .C(
        \counter[4]_net_1 ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] ));
    NOR2A \off_reg_RNI3C43[4]  (.A(\off_reg[4]_net_1 ), .B(act_ctl_5_2)
        , .Y(\off_time[4] ));
    NOR2A \counter_RNO_1[31]  (.A(\counter[31]_net_1 ), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(N_322));
    OR2B un1_counter_2_0_I_133 (.A(N_2), .B(\counter[2]_net_1 ), .Y(
        N_8));
    DFN1C0 \counter[14]  (.D(counter_n14), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[14]_net_1 ));
    DFN1E1C0 \off_reg[29]  (.D(off_div[29]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[29]_net_1 ));
    AND3 un1_counter_2_0_I_18 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[0] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] ));
    DFN1E1C0 \off_reg[1]  (.D(off_div[1]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[1]_net_1 ));
    NOR2A \off_reg_RNIOETI[22]  (.A(\off_reg[22]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[22] ));
    NOR2A \counter_RNO[22]  (.A(counter_n22_tz), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n22));
    NOR3C \counter_RNIL7BH4[10]  (.A(\counter[9]_net_1 ), .B(
        counter_c8), .C(\counter[10]_net_1 ), .Y(counter_c10));
    AO1C un1_counter_0_I_131 (.A(\off_time[1] ), .B(\counter[1]_net_1 )
        , .C(N_4_0), .Y(N_6_0));
    AND2 un1_counter_0_I_19 (.A(\DWACT_BL_EQUAL_0_E[12] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[3] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[1] ));
    NOR2B \counter_RNICOCS4[11]  (.A(counter_c10), .B(
        \counter[11]_net_1 ), .Y(counter_c11));
    XNOR2 un1_counter_0_I_42 (.A(\counter[26]_net_1 ), .B(
        \off_time[26] ), .Y(\DWACT_BL_EQUAL_0_E_3[2] ));
    AO1C un1_counter_0_I_135 (.A(\counter[3]_net_1 ), .B(\off_time[3] )
        , .C(N_5), .Y(N_10_0));
    DFN1E1C0 \off_reg[10]  (.D(off_div[10]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[10]_net_1 ));
    NOR2A un1_counter_0_I_85 (.A(\off_time[15] ), .B(
        \counter[15]_net_1 ), .Y(\ACT_LT4_E[0] ));
    DFN1C0 \counter[31]  (.D(counter_n31), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[31]_net_1 ));
    OR2A un1_counter_0_I_32 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .Y(N_43));
    OA1A un1_counter_0_I_62 (.A(N_36), .B(N_38), .C(N_37), .Y(N_41));
    OA1 un1_counter_0_I_137 (.A(N_11_0), .B(N_10_0), .C(N_9), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] ));
    AO1 un1_counter_0_I_138 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_1[2] ));
    NOR2A \off_reg_RNINDTI[21]  (.A(\off_reg[21]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[21] ));
    NOR2A \off_reg_RNI0943[1]  (.A(\off_reg[1]_net_1 ), .B(act_ctl_5_2)
        , .Y(\off_time[1] ));
    NOR3C \counter_RNIVKSV7[19]  (.A(\counter[19]_net_1 ), .B(
        counter_c18), .C(\counter[20]_net_1 ), .Y(counter_c20));
    NOR2A un1_counter_0_I_92 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\ACT_LT4_E[7] ));
    OR2 \off_reg_RNI9K74[9]  (.A(\off_reg[9]_net_1 ), .B(act_ctl_5_3), 
        .Y(\off_time[9] ));
    DFN1C0 \counter[24]  (.D(counter_n24), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[24]_net_1 ));
    OR2A un1_counter_0_I_119 (.A(\off_time[9] ), .B(\counter[9]_net_1 )
        , .Y(N_15));
    NOR3 un1_counter_2_0_I_14 (.A(\counter[29]_net_1 ), .B(
        \counter[30]_net_1 ), .C(\counter[28]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[3] ));
    AND3 un1_counter_2_0_I_78 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ));
    NOR2B \counter_RNIR2L3B[29]  (.A(counter_c28), .B(
        \counter[29]_net_1 ), .Y(counter_c29));
    XNOR2 un1_counter_0_I_80 (.A(\counter[17]_net_1 ), .B(
        \off_time[17] ), .Y(\DWACT_BL_EQUAL_0_E_1[2] ));
    XNOR2 un1_counter_0_I_5 (.A(\counter[27]_net_1 ), .B(
        \off_time[27] ), .Y(\DWACT_BL_EQUAL_0_E_0[8] ));
    AND3 un1_counter_0_I_113 (.A(\DWACT_BL_EQUAL_0_E_0[0] ), .B(
        \DWACT_BL_EQUAL_0_E_0[1] ), .C(\DWACT_BL_EQUAL_0_E_0[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] ));
    XNOR2 un1_counter_0_I_24 (.A(\counter[28]_net_1 ), .B(
        \off_time[28] ), .Y(\DWACT_BL_EQUAL_0_E_4[1] ));
    NOR2A \counter_RNO[4]  (.A(counter_n4_tz), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n4));
    AND3 un1_counter_0_I_75 (.A(\DWACT_BL_EQUAL_0_E[6] ), .B(
        \DWACT_BL_EQUAL_0_E[7] ), .C(\DWACT_BL_EQUAL_0_E[8] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[2] ));
    DFN1E1C0 \off_reg[14]  (.D(off_div[14]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[14]_net_1 ));
    NOR3C \counter_RNIAIE33[11]  (.A(counter_m6_0_a2_2), .B(
        counter_m6_0_a2_1), .C(counter_m6_0_a2_6), .Y(
        counter_m6_0_a2_7));
    AO1B un1_counter_2_0_I_120 (.A(act_ctl_5_0), .B(\counter[6]_net_1 )
        , .C(N_14), .Y(N_16));
    XA1B \counter_RNO[18]  (.A(\counter[18]_net_1 ), .B(counter_c17), 
        .C(N_403_0), .Y(counter_n18));
    NOR3 un1_counter_2_0_I_15 (.A(\counter[26]_net_1 ), .B(
        \counter[27]_net_1 ), .C(\counter[25]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[2] ));
    OR2A un1_counter_0_I_86 (.A(\off_time[16] ), .B(
        \counter[16]_net_1 ), .Y(\ACT_LT4_E[1] ));
    OA1A un1_counter_0_I_58 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .C(N_33), .Y(N_37));
    OA1A un1_counter_0_I_121 (.A(\counter[8]_net_1 ), .B(\off_time[8] )
        , .C(N_13_0), .Y(N_17_0));
    OR2 \off_reg_RNITISI[18]  (.A(\off_reg[18]_net_1 ), .B(act_ctl_5_7)
        , .Y(\off_time[18] ));
    AND2 un1_counter_2_0_I_20 (.A(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[1] ), .B(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E[0] ), .Y(
        \DWACT_COMP0_E[1] ));
    AX1C \counter_RNO_0[26]  (.A(\counter[25]_net_1 ), .B(counter_c24), 
        .C(\counter[26]_net_1 ), .Y(counter_n26_tz));
    XA1B \counter_RNO[27]  (.A(\counter[27]_net_1 ), .B(counter_c26), 
        .C(N_403_0), .Y(counter_n27));
    OA1A un1_counter_0_I_125 (.A(N_16_0), .B(N_18_0), .C(N_17_0), .Y(
        N_21_0));
    AX1C \counter_RNO_0[6]  (.A(\counter[5]_net_1 ), .B(counter_c4), 
        .C(\counter[6]_net_1 ), .Y(counter_n6_tz));
    XNOR2 un1_counter_0_I_70 (.A(\counter[15]_net_1 ), .B(
        \off_time[15] ), .Y(\DWACT_BL_EQUAL_0_E[5] ));
    OA1 un1_counter_0_I_106 (.A(N_31), .B(N_30), .C(N_29), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] ));
    DFN1E1C0 \off_reg[18]  (.D(off_div[18]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[18]_net_1 ));
    AO1C un1_counter_0_I_102 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .C(N_22), .Y(N_28));
    OR2B un1_counter_2_0_I_117 (.A(act_ctl_5_3), .B(\counter[7]_net_1 )
        , .Y(N_13));
    AND3 un1_counter_2_0_I_113 (.A(\DWACT_BL_EQUAL_0_E[0] ), .B(
        \DWACT_BL_EQUAL_0_E[1] ), .C(\DWACT_BL_EQUAL_0_E[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ));
    XNOR2 un1_counter_0_I_44 (.A(\counter[24]_net_1 ), .B(
        \off_time[24] ), .Y(\DWACT_BL_EQUAL_0_E_3[0] ));
    OR2A un1_counter_0_I_53 (.A(\off_time[20] ), .B(
        \counter[20]_net_1 ), .Y(N_32));
    OR2A un1_counter_0_I_127 (.A(\off_time[1] ), .B(\counter[1]_net_1 )
        , .Y(N_2_0));
    OR2A un1_counter_0_I_34 (.A(\off_time[31] ), .B(
        \counter[31]_net_1 ), .Y(N_45));
    OR2A un1_counter_0_I_128 (.A(\counter[2]_net_1 ), .B(\off_time[2] )
        , .Y(N_3));
    OR2A un1_counter_0_I_89 (.A(\off_time[17] ), .B(
        \counter[17]_net_1 ), .Y(\ACT_LT4_E[4] ));
    AO1 un1_counter_0_I_64 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_3[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_3[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[2] ));
    DFN1E1C0 \off_reg[16]  (.D(off_div[16]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[16]_net_1 ));
    AND3 un1_counter_0_I_76 (.A(\DWACT_BL_EQUAL_0_E_1[3] ), .B(
        \DWACT_BL_EQUAL_0_E_0[4] ), .C(\DWACT_BL_EQUAL_0_E[5] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[1] ));
    XNOR2 un1_counter_0_I_1 (.A(\counter[23]_net_1 ), .B(
        \off_time[23] ), .Y(\DWACT_BL_EQUAL_0_E_2[4] ));
    DFN1E1C0 \off_reg[30]  (.D(off_div[30]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[30]_net_1 ));
    NOR3C \counter_RNIHQRO3[8]  (.A(\counter[7]_net_1 ), .B(counter_c6)
        , .C(\counter[8]_net_1 ), .Y(counter_c8));
    NOR3 un1_counter_2_0_I_75 (.A(\counter[17]_net_1 ), .B(
        \counter[18]_net_1 ), .C(\counter[16]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[2] ));
    NOR2A \off_reg_RNIPI1K[31]  (.A(\off_reg[31]_net_1 ), .B(
        act_ctl_5_8), .Y(\off_time[31] ));
    NOR2A \counter_RNO[24]  (.A(counter_n24_tz), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n24));
    DFN1C0 \counter[7]  (.D(counter_n7), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[7]_net_1 ));
    AOI1A un1_counter_0_I_94 (.A(\ACT_LT4_E[7] ), .B(\ACT_LT4_E[8] ), 
        .C(\ACT_LT4_E[5] ), .Y(\ACT_LT4_E[10] ));
    DFN1C0 \counter[30]  (.D(counter_n30), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[30]_net_1 ));
    NOR2A \off_reg_RNINCSI[12]  (.A(\off_reg[12]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[12] ));
    OA1 un1_counter_0_I_41 (.A(N_51), .B(N_50), .C(N_49), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E_0[0] ));
    AND3 un1_counter_0_I_18 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_6[0] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_5[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[2] ), .Y(
        \DWACT_BL_ANDTREE_0_DWACT_BL_ANDTREE_0_E_0[0] ));
    NOR2B \counter_RNI4AE75[12]  (.A(counter_c11), .B(
        \counter[12]_net_1 ), .Y(counter_c12));
    OR2A un1_counter_0_I_31 (.A(\off_time[28] ), .B(
        \counter[28]_net_1 ), .Y(N_42));
    NOR2A \off_reg_RNIV743[0]  (.A(\off_reg[0]_net_1 ), .B(act_ctl_5_2)
        , .Y(\off_time[0] ));
    NOR3C \counter_RNI567C9[24]  (.A(\counter[23]_net_1 ), .B(
        counter_c22), .C(\counter[24]_net_1 ), .Y(counter_c24));
    XNOR2 un1_counter_2_0_I_108 (.A(\counter[5]_net_1 ), .B(
        act_ctl_5_3), .Y(\DWACT_BL_EQUAL_0_E[0] ));
    AO1C un1_counter_0_I_61 (.A(\counter[22]_net_1 ), .B(
        \off_time[22] ), .C(N_35), .Y(N_40));
    NOR2 \counter_RNO[0]  (.A(\counter[0]_net_1 ), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(\counter_RNO_3[0] ));
    XNOR2 un1_counter_0_I_79 (.A(\counter[18]_net_1 ), .B(
        \off_time[18] ), .Y(\DWACT_BL_EQUAL_0_E_0[3] ));
    DFN1E1C0 \off_reg[3]  (.D(off_div[3]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[3]_net_1 ));
    DFN1E1C0 \off_reg[0]  (.D(off_div[0]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[0]_net_1 ));
    NOR2A un1_counter_2_0_I_126 (.A(N_21), .B(\counter[9]_net_1 ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ));
    OR2A un1_counter_0_I_134 (.A(\counter[4]_net_1 ), .B(\off_time[4] )
        , .Y(N_9));
    XNOR2 un1_counter_0_I_13 (.A(\counter[28]_net_1 ), .B(
        \off_time[28] ), .Y(\DWACT_BL_EQUAL_0_E[9] ));
    NOR2A un1_counter_0_I_91 (.A(\ACT_LT4_E[4] ), .B(\ACT_LT4_E[5] ), 
        .Y(\ACT_LT4_E[6] ));
    NOR2A \off_reg_RNI1A43[2]  (.A(\off_reg[2]_net_1 ), .B(act_ctl_5_2)
        , .Y(\off_time[2] ));
    AOI1A un1_counter_0_I_52 (.A(\ACT_LT3_E[3] ), .B(\ACT_LT3_E[4] ), 
        .C(\ACT_LT3_E[5] ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E_2[0] ));
    NOR2A \counter_RNO[20]  (.A(counter_n20_tz), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n20));
    NOR2A \off_reg_RNIMBSI[11]  (.A(\off_reg[11]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[11] ));
    OR2 \off_reg_RNI5E43[6]  (.A(\off_reg[6]_net_1 ), .B(act_ctl_5_2), 
        .Y(\off_time[6] ));
    DFN1E1C0 \off_reg[13]  (.D(off_div[13]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[13]_net_1 ));
    XNOR2 un1_counter_0_I_27 (.A(\counter[31]_net_1 ), .B(
        \off_time[31] ), .Y(\DWACT_BL_EQUAL_0_E_1[4] ));
    XNOR2 un1_counter_0_I_111 (.A(\counter[7]_net_1 ), .B(
        \off_time[7] ), .Y(\DWACT_BL_EQUAL_0_E_0[2] ));
    OA1A un1_counter_2_0_I_136 (.A(N_6), .B(N_8), .C(N_7), .Y(N_11));
    AND2 un1_counter_0_I_115 (.A(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[1] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_2[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E_2[1] ));
    DFN1E1C0 \off_reg[4]  (.D(off_div[4]), .CLK(clk_c), .CLR(n_rst_c), 
        .E(pwm_chg_0), .Q(\off_reg[4]_net_1 ));
    XNOR2 un1_counter_0_I_8 (.A(\counter[25]_net_1 ), .B(
        \off_time[25] ), .Y(\DWACT_BL_EQUAL_0_E_0[6] ));
    DFN1E1C0 \off_reg[20]  (.D(off_div[20]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[20]_net_1 ));
    NOR2A \counter_RNO[2]  (.A(counter_n2_tz), .B(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n2));
    NOR3C \counter_RNIUKC2A[26]  (.A(\counter[25]_net_1 ), .B(
        counter_c24), .C(\counter[26]_net_1 ), .Y(counter_c26));
    DFN1C0 \counter[9]  (.D(counter_n9), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[9]_net_1 ));
    NOR3 un1_counter_2_0_I_16 (.A(\counter[24]_net_1 ), .B(
        \counter[23]_net_1 ), .C(\counter[22]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_1[1] ));
    NOR2 un1_counter_2_0_I_114 (.A(\counter[8]_net_1 ), .B(
        \counter[9]_net_1 ), .Y(\DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ));
    OR2A un1_counter_0_I_117 (.A(\counter[7]_net_1 ), .B(\off_time[7] )
        , .Y(N_13_0));
    XA1B \counter_RNO[19]  (.A(\counter[19]_net_1 ), .B(counter_c18), 
        .C(N_403_0), .Y(counter_n19));
    AO1C un1_counter_0_I_124 (.A(\counter[8]_net_1 ), .B(\off_time[8] )
        , .C(N_15), .Y(N_20));
    NOR2A un1_counter_0_I_118 (.A(\off_time[5] ), .B(
        \counter[5]_net_1 ), .Y(N_14_0));
    XNOR2 un1_counter_0_I_12 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .Y(\DWACT_BL_EQUAL_0_E_5[2] ));
    AO1 un1_counter_2_0_I_138 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[1] )
        , .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E_0[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] ));
    NOR2A \off_reg_RNI2B43[3]  (.A(\off_reg[3]_net_1 ), .B(act_ctl_5_2)
        , .Y(\off_time[3] ));
    XA1B \counter_RNO[9]  (.A(\counter[9]_net_1 ), .B(counter_c8), .C(
        cur_pwm_RNI9RT933_0_net_1), .Y(counter_n9));
    NOR2B \counter_RNII5J86[15]  (.A(counter_c14), .B(
        \counter[15]_net_1 ), .Y(counter_c15));
    DFN1E1C0 \off_reg[12]  (.D(off_div[12]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg_0), .Q(\off_reg[12]_net_1 ));
    AOI1A un1_counter_0_I_88 (.A(\ACT_LT4_E[0] ), .B(\ACT_LT4_E[1] ), 
        .C(\ACT_LT4_E[2] ), .Y(\ACT_LT4_E[3] ));
    OR2A un1_counter_0_I_47 (.A(\off_time[25] ), .B(
        \counter[25]_net_1 ), .Y(\ACT_LT3_E[1] ));
    DFN1C0 \counter[8]  (.D(counter_n8), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[8]_net_1 ));
    NOR2A \off_reg_RNIVN0K[28]  (.A(\off_reg[28]_net_1 ), .B(
        act_ctl_5_8), .Y(\off_time[28] ));
    OR2A un1_counter_0_I_54 (.A(\counter[21]_net_1 ), .B(
        \off_time[21] ), .Y(N_33));
    AO1C un1_counter_0_I_37 (.A(\counter[29]_net_1 ), .B(
        \off_time[29] ), .C(N_42), .Y(N_48));
    OR2 \off_reg_RNIUJSI[19]  (.A(\off_reg[19]_net_1 ), .B(act_ctl_5_7)
        , .Y(\off_time[19] ));
    NOR2A \off_reg_RNIQFSI[15]  (.A(\off_reg[15]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[15] ));
    XNOR2 un1_counter_0_I_7 (.A(\counter[26]_net_1 ), .B(
        \off_time[26] ), .Y(\DWACT_BL_EQUAL_0_E_0[7] ));
    XNOR2 un1_counter_0_I_67 (.A(\counter[14]_net_1 ), .B(
        \off_time[14] ), .Y(\DWACT_BL_EQUAL_0_E_0[4] ));
    DFN1C0 \counter[18]  (.D(counter_n18), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\counter[18]_net_1 ));
    AO1C un1_counter_0_I_100 (.A(\off_time[11] ), .B(
        \counter[11]_net_1 ), .C(N_24), .Y(N_26));
    DFN1E1C0 \off_reg[24]  (.D(off_div[24]), .CLK(clk_c), .CLR(n_rst_c)
        , .E(pwm_chg), .Q(\off_reg[24]_net_1 ));
    AND3 un1_counter_0_I_83 (.A(\DWACT_BL_EQUAL_0_E_1[0] ), .B(
        \DWACT_BL_EQUAL_0_E_1[1] ), .C(\DWACT_BL_EQUAL_0_E_1[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_3[0] ));
    MX2C cur_pwm_RNI9RT933 (.A(I_140_8), .B(I_140_7), .S(primary_15_c), 
        .Y(N_403_0));
    XA1B \counter_RNO[16]  (.A(\counter[16]_net_1 ), .B(counter_c15), 
        .C(N_403_0), .Y(counter_n16));
    DFN1C0 \counter[0]  (.D(\counter_RNO_3[0] ), .CLK(clk_c), .CLR(
        n_rst_c), .Q(\counter[0]_net_1 ));
    NOR3 un1_counter_2_0_I_76 (.A(\counter[15]_net_1 ), .B(
        \counter[14]_net_1 ), .C(\counter[13]_net_1 ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[1] ));
    OR2A un1_counter_0_I_97 (.A(\counter[12]_net_1 ), .B(
        \off_time[12] ), .Y(N_23));
    NOR2A \off_reg_RNISK0K[25]  (.A(\off_reg[25]_net_1 ), .B(
        act_ctl_5_8), .Y(\off_time[25] ));
    NOR2A \off_reg_RNIPFTI[23]  (.A(\off_reg[23]_net_1 ), .B(
        act_ctl_5_7), .Y(\off_time[23] ));
    
endmodule


module spi_clk_11s_3_1(
       sck_5_c,
       n_rst_c,
       clk_c
    );
output sck_5_c;
input  n_rst_c;
input  clk_c;

    wire N_8, \counter[1]_net_1 , \counter[0]_net_1 , N_6, 
        \counter[3]_net_1 , \DWACT_FINC_E[0] , cur_clk5_5, cur_clk5_3, 
        \counter[6]_net_1 , cur_clk5_4, cur_clk5_1, \counter[7]_net_1 , 
        \counter[8]_net_1 , \counter[4]_net_1 , \counter[5]_net_1 , 
        \counter[2]_net_1 , cur_clk_RNO_3, \counter_3[1] , I_5_3, 
        \counter_3[0] , \counter_3[3] , I_9_3, I_7_3, I_12_4, I_14_7, 
        I_17_4, I_20_7, I_23_10, N_2, \DWACT_FINC_E[2] , 
        \DWACT_FINC_E[3] , N_3, N_4, \DWACT_FINC_E[1] , N_5, N_7, GND, 
        VCC;
    
    NOR2B un3_counter_I_6 (.A(\counter[1]_net_1 ), .B(
        \counter[0]_net_1 ), .Y(N_8));
    AND3 un3_counter_I_19 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\counter[6]_net_1 ), .Y(N_3));
    XOR2 un3_counter_I_20 (.A(N_3), .B(\counter[7]_net_1 ), .Y(I_20_7));
    DFN1C0 \counter[2]  (.D(I_7_3), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[2]_net_1 ));
    DFN1C0 \counter[7]  (.D(I_20_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[7]_net_1 ));
    AND3 un3_counter_I_13 (.A(\DWACT_FINC_E[0] ), .B(
        \counter[3]_net_1 ), .C(\counter[4]_net_1 ), .Y(N_5));
    NOR3A \counter_RNI6G52[8]  (.A(cur_clk5_1), .B(\counter[7]_net_1 ), 
        .C(\counter[8]_net_1 ), .Y(cur_clk5_4));
    AOI1 \counter_RNO[0]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(
        \counter[0]_net_1 ), .Y(\counter_3[0] ));
    DFN1C0 \counter[6]  (.D(I_17_4), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[6]_net_1 ));
    VCC VCC_i (.Y(VCC));
    XOR2 un3_counter_I_12 (.A(N_6), .B(\counter[4]_net_1 ), .Y(I_12_4));
    DFN1C0 \counter[8]  (.D(I_23_10), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[8]_net_1 ));
    XOR2 un3_counter_I_23 (.A(N_2), .B(\counter[8]_net_1 ), .Y(I_23_10)
        );
    AOI1B \counter_RNO[1]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(I_5_3), 
        .Y(\counter_3[1] ));
    AND3 un3_counter_I_22 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[2] )
        , .C(\DWACT_FINC_E[3] ), .Y(N_2));
    XOR2 un3_counter_I_7 (.A(N_8), .B(\counter[2]_net_1 ), .Y(I_7_3));
    NOR2B un3_counter_I_11 (.A(\counter[3]_net_1 ), .B(
        \DWACT_FINC_E[0] ), .Y(N_6));
    AND3 un3_counter_I_16 (.A(\DWACT_FINC_E[0] ), .B(\DWACT_FINC_E[1] )
        , .C(\counter[5]_net_1 ), .Y(N_4));
    DFN1C0 \counter[4]  (.D(I_12_4), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[4]_net_1 ));
    XOR2 un3_counter_I_17 (.A(N_4), .B(\counter[6]_net_1 ), .Y(I_17_4));
    NOR2A \counter_RNIVJ21[4]  (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(cur_clk5_3));
    DFN1C0 \counter[5]  (.D(I_14_7), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \counter[5]_net_1 ));
    AND3 un3_counter_I_8 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(N_7));
    GND GND_i (.Y(GND));
    AX1C cur_clk_RNO (.A(cur_clk5_4), .B(cur_clk5_5), .C(sck_5_c), .Y(
        cur_clk_RNO_3));
    AOI1B \counter_RNO[3]  (.A(cur_clk5_5), .B(cur_clk5_4), .C(I_9_3), 
        .Y(\counter_3[3] ));
    AND2 un3_counter_I_21 (.A(\counter[6]_net_1 ), .B(
        \counter[7]_net_1 ), .Y(\DWACT_FINC_E[3] ));
    DFN1C0 \counter[1]  (.D(\counter_3[1] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[1]_net_1 ));
    DFN1C0 \counter[3]  (.D(\counter_3[3] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[3]_net_1 ));
    NOR2 \counter_RNIVJ21[2]  (.A(\counter[5]_net_1 ), .B(
        \counter[2]_net_1 ), .Y(cur_clk5_1));
    NOR3B \counter_RNIU752[6]  (.A(\counter[1]_net_1 ), .B(cur_clk5_3), 
        .C(\counter[6]_net_1 ), .Y(cur_clk5_5));
    AND2 un3_counter_I_15 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .Y(\DWACT_FINC_E[1] ));
    XOR2 un3_counter_I_9 (.A(N_7), .B(\counter[3]_net_1 ), .Y(I_9_3));
    DFN1C0 cur_clk (.D(cur_clk_RNO_3), .CLK(clk_c), .CLR(n_rst_c), .Q(
        sck_5_c));
    XOR2 un3_counter_I_14 (.A(N_5), .B(\counter[5]_net_1 ), .Y(I_14_7));
    XOR2 un3_counter_I_5 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .Y(I_5_3));
    AND3 un3_counter_I_10 (.A(\counter[0]_net_1 ), .B(
        \counter[1]_net_1 ), .C(\counter[2]_net_1 ), .Y(
        \DWACT_FINC_E[0] ));
    DFN1C0 \counter[0]  (.D(\counter_3[0] ), .CLK(clk_c), .CLR(n_rst_c)
        , .Q(\counter[0]_net_1 ));
    AND3 un3_counter_I_18 (.A(\counter[3]_net_1 ), .B(
        \counter[4]_net_1 ), .C(\counter[5]_net_1 ), .Y(
        \DWACT_FINC_E[2] ));
    
endmodule


module PID_controller_Z5(
       LED_15,
       primary_15_c,
       act_ctl_5_3,
       act_ctl_5_4,
       act_ctl_5_2,
       act_ctl_5_7,
       act_ctl_5_8,
       act_ctl_5_0,
       din_15_c,
       cs_i_1_i,
       sck_5_c,
       clk_c,
       n_rst_c
    );
output [7:0] LED_15;
output primary_15_c;
input  act_ctl_5_3;
input  act_ctl_5_4;
input  act_ctl_5_2;
input  act_ctl_5_7;
input  act_ctl_5_8;
input  act_ctl_5_0;
input  din_15_c;
output cs_i_1_i;
output sck_5_c;
input  clk_c;
input  n_rst_c;

    wire pwm_chg, N_46_1, N_46_1_0, sig_prev, sig_old_i_0, pwm_rdy, 
        sig_old_i_0_0, sig_prev_0, sum_rdy, deriv_enable, calc_avg, 
        calc_int, pwm_enable, sum_enable, calc_error, avg_enable, 
        int_enable, pwm_chg_0, avg_enable_0, avg_enable_1, \cur_vd[0] , 
        \cur_vd[1] , \cur_vd[2] , \cur_vd[3] , \cur_vd[4] , 
        \cur_vd[5] , \cur_vd[6] , \cur_vd[7] , \cur_vd[8] , 
        \cur_vd[9] , \cur_vd[10] , \cur_vd[11] , \avg_new[0] , 
        \avg_new[1] , \avg_new[2] , \avg_new[3] , \avg_new[4] , 
        \avg_new[5] , \avg_new[6] , \avg_new[7] , \avg_new[8] , 
        \avg_new[9] , \avg_new[10] , \avg_new[11] , \avg_old[0] , 
        \avg_old[1] , \avg_old[2] , \avg_old[3] , \avg_old[4] , 
        \avg_old[5] , \avg_old[6] , \avg_old[7] , \avg_old[8] , 
        \avg_old[9] , \avg_old[10] , \avg_old[11] , \cur_error[0] , 
        \cur_error[1] , \cur_error[2] , \cur_error[3] , \cur_error[4] , 
        \cur_error[5] , \cur_error[6] , \cur_error[7] , \cur_error[8] , 
        \cur_error[9] , \cur_error[10] , \cur_error[11] , 
        \cur_error[12] , \LED_15_i[5] , \average[2] , \average[3] , 
        \average[4] , \average[5] , \average[6] , \sr_old[0] , 
        \sr_old[1] , \sr_old[2] , \sr_old[3] , \sr_old[4] , 
        \sr_old[5] , \sr_old[6] , \sr_old[7] , \sr_old[8] , 
        \sr_old[9] , \sr_old[10] , \sr_old[11] , \sr_old[12] , 
        \sr_new[0] , \sr_new[1] , \sr_new[2] , \sr_new[3] , 
        \sr_new[4] , \sr_new[5] , \sr_new[6] , \sr_new[7] , 
        \sr_new[8] , \sr_new[9] , \sr_new[10] , \sr_new[11] , 
        \sr_new[12] , \sr_prev[0] , \sr_prev[1] , \sr_prev[2] , 
        \sr_prev[3] , \sr_prev[4] , \sr_prev[5] , \sr_prev[6] , 
        \sr_prev[7] , \sr_prev[8] , \sr_prev[9] , \sr_prev[10] , 
        \sr_prev[11] , \sr_prev[12] , \sr_new_0[12] , \integral[6] , 
        \integral[7] , \integral[8] , \integral[9] , \integral[10] , 
        \integral[11] , \integral[12] , \integral[13] , \integral[14] , 
        \integral[15] , \integral[16] , \integral[17] , \integral[18] , 
        \integral[19] , \integral[20] , \integral[21] , \integral[22] , 
        \integral[23] , \integral[24] , \integral[25] , 
        \integral_i[24] , \integral_i[25] , \integral_0[25] , 
        \integral_1[25] , \derivative[12] , \sum[39] , \sum[14] , 
        \sum[20] , \sum[19] , \sum[22] , \sum[13] , \sum[17] , 
        \sum[18] , \sum[23] , \sum[21] , \sum[16] , \sum[15] , 
        \sum[12] , \sum[11] , \sum[6] , \sum[9] , \sum[10] , \sum[5] , 
        \sum[8] , \sum[7] , \sum[4] , \sum[2] , \sum[1] , \sum[0] , 
        \sum[3] , \sum_0[39] , \sum_1[39] , \sum_2[39] , vd_done, 
        \off_div[0] , \off_div[1] , \off_div[2] , \off_div[3] , 
        \off_div[4] , \off_div[5] , \off_div[6] , \off_div[7] , 
        \off_div[8] , \off_div[9] , \off_div[10] , \off_div[11] , 
        \off_div[12] , \off_div[13] , \off_div[14] , \off_div[15] , 
        \off_div[16] , \off_div[17] , \off_div[18] , \off_div[19] , 
        \off_div[20] , \off_div[21] , \off_div[22] , \off_div[23] , 
        \off_div[24] , \off_div[25] , \off_div[26] , \off_div[27] , 
        \off_div[28] , \off_div[29] , \off_div[30] , \off_div[31] , 
        GND, VCC;
    
    pwm_ctl_200s_32s_13s_0_1_2_2 PWM_CTL (.sum_8(\sum[8] ), .sum_39(
        \sum[39] ), .sum_10(\sum[10] ), .sum_11(\sum[11] ), .sum_12(
        \sum[12] ), .sum_13(\sum[13] ), .sum_15(\sum[15] ), .sum_16(
        \sum[16] ), .sum_17(\sum[17] ), .sum_18(\sum[18] ), .sum_19(
        \sum[19] ), .sum_20(\sum[20] ), .sum_21(\sum[21] ), .sum_22(
        \sum[22] ), .sum_23(\sum[23] ), .sum_14(\sum[14] ), .sum_9(
        \sum[9] ), .sum_2_d0(\sum[2] ), .sum_1_d0(\sum[1] ), .sum_0_d0(
        \sum[0] ), .sum_7(\sum[7] ), .sum_6(\sum[6] ), .sum_4(\sum[4] )
        , .sum_3(\sum[3] ), .sum_5(\sum[5] ), .off_div({\off_div[31] , 
        \off_div[30] , \off_div[29] , \off_div[28] , \off_div[27] , 
        \off_div[26] , \off_div[25] , \off_div[24] , \off_div[23] , 
        \off_div[22] , \off_div[21] , \off_div[20] , \off_div[19] , 
        \off_div[18] , \off_div[17] , \off_div[16] , \off_div[15] , 
        \off_div[14] , \off_div[13] , \off_div[12] , \off_div[11] , 
        \off_div[10] , \off_div[9] , \off_div[8] , \off_div[7] , 
        \off_div[6] , \off_div[5] , \off_div[4] , \off_div[3] , 
        \off_div[2] , \off_div[1] , \off_div[0] }), .sum_1_0(
        \sum_1[39] ), .sum_0_0(\sum_0[39] ), .sum_2_0(\sum_2[39] ), 
        .n_rst_c(n_rst_c), .clk_c(clk_c), .pwm_enable(pwm_enable), 
        .pwm_rdy(pwm_rdy));
    integral_calc_13s_4_3 AVG_CALC (.avg_old({\avg_old[11] , 
        \avg_old[10] , \avg_old[9] , \avg_old[8] , \avg_old[7] , 
        \avg_old[6] , \avg_old[5] , \avg_old[4] , \avg_old[3] , 
        \avg_old[2] , \avg_old[1] , \avg_old[0] }), .avg_new({
        \avg_new[11] , \avg_new[10] , \avg_new[9] , \avg_new[8] , 
        \avg_new[7] , \avg_new[6] , \avg_new[5] , \avg_new[4] , 
        \avg_new[3] , \avg_new[2] , \avg_new[1] , \avg_new[0] }), 
        .average({\average[6] , \average[5] , \average[4] , 
        \average[3] , \average[2] }), .LED_15({LED_15[7], LED_15[6], 
        LED_15[5], LED_15[4], LED_15[3], LED_15[2], LED_15[1], 
        LED_15[0]}), .LED_15_i_0(\LED_15_i[5] ), .calc_avg(calc_avg), 
        .N_46_1(N_46_1), .n_rst_c(n_rst_c), .clk_c(clk_c));
    error_sr_13s_5s_3 AVGSR (.cur_vd({\cur_vd[11] , \cur_vd[10] , 
        \cur_vd[9] , \cur_vd[8] , \cur_vd[7] , \cur_vd[6] , 
        \cur_vd[5] , \cur_vd[4] , \cur_vd[3] , \cur_vd[2] , 
        \cur_vd[1] , \cur_vd[0] }), .avg_new({\avg_new[11] , 
        \avg_new[10] , \avg_new[9] , \avg_new[8] , \avg_new[7] , 
        \avg_new[6] , \avg_new[5] , \avg_new[4] , \avg_new[3] , 
        \avg_new[2] , \avg_new[1] , \avg_new[0] }), .avg_old({
        \avg_old[11] , \avg_old[10] , \avg_old[9] , \avg_old[8] , 
        \avg_old[7] , \avg_old[6] , \avg_old[5] , \avg_old[4] , 
        \avg_old[3] , \avg_old[2] , \avg_old[1] , \avg_old[0] }), 
        .avg_enable_0(avg_enable_0), .avg_enable(avg_enable), 
        .avg_enable_1(avg_enable_1), .n_rst_c(n_rst_c), .clk_c(clk_c));
    error_sr_13s_64s_3 INTSR (.sr_old({\sr_old[12] , \sr_old[11] , 
        \sr_old[10] , \sr_old[9] , \sr_old[8] , \sr_old[7] , 
        \sr_old[6] , \sr_old[5] , \sr_old[4] , \sr_old[3] , 
        \sr_old[2] , \sr_old[1] , \sr_old[0] }), .sr_new({\sr_new[12] , 
        \sr_new[11] , \sr_new[10] , \sr_new[9] , \sr_new[8] , 
        \sr_new[7] , \sr_new[6] , \sr_new[5] , \sr_new[4] , 
        \sr_new[3] , \sr_new[2] , \sr_new[1] , \sr_new[0] }), 
        .cur_error({\cur_error[12] , \cur_error[11] , \cur_error[10] , 
        \cur_error[9] , \cur_error[8] , \cur_error[7] , \cur_error[6] , 
        \cur_error[5] , \cur_error[4] , \cur_error[3] , \cur_error[2] , 
        \cur_error[1] , \cur_error[0] }), .sr_prev({\sr_prev[12] , 
        \sr_prev[11] , \sr_prev[10] , \sr_prev[9] , \sr_prev[8] , 
        \sr_prev[7] , \sr_prev[6] , \sr_prev[5] , \sr_prev[4] , 
        \sr_prev[3] , \sr_prev[2] , \sr_prev[1] , \sr_prev[0] }), 
        .sr_new_0_0(\sr_new_0[12] ), .int_enable(int_enable), .n_rst_c(
        n_rst_c), .clk_c(clk_c));
    controller_Z1_4_3 CONTROLLER (.pwm_chg(pwm_chg), .N_46_1_0(N_46_1), 
        .N_46_1(N_46_1_0), .sig_prev_0(sig_prev), .sig_old_i_0_0(
        sig_old_i_0), .pwm_rdy(pwm_rdy), .sig_old_i_0(sig_old_i_0_0), 
        .sig_prev(sig_prev_0), .sum_rdy(sum_rdy), .deriv_enable(
        deriv_enable), .calc_avg(calc_avg), .calc_int(calc_int), 
        .pwm_enable(pwm_enable), .sum_enable(sum_enable), .calc_error(
        calc_error), .avg_enable(avg_enable), .int_enable(int_enable), 
        .pwm_chg_0(pwm_chg_0), .avg_enable_0(avg_enable_0), .n_rst_c(
        n_rst_c), .clk_c(clk_c), .avg_enable_1(avg_enable_1));
    sig_gen_8 FM_CYCLE (.primary_15_c(primary_15_c), .n_rst_c(n_rst_c), 
        .clk_c(clk_c), .sig_old_i_0(sig_old_i_0), .sig_prev(sig_prev));
    pid_sum_13s_4_3 SUM (.integral_i({\integral_i[25] , 
        \integral_i[24] }), .integral({\integral[25] , \integral[24] , 
        \integral[23] , \integral[22] , \integral[21] , \integral[20] , 
        \integral[19] , \integral[18] , \integral[17] , \integral[16] , 
        \integral[15] , \integral[14] , \integral[13] , \integral[12] , 
        \integral[11] , \integral[10] , \integral[9] , \integral[8] , 
        \integral[7] , \integral[6] }), .derivative_0(\derivative[12] )
        , .sr_new({\sr_new[12] , \sr_new[11] , \sr_new[10] , 
        \sr_new[9] , \sr_new[8] , \sr_new[7] , \sr_new[6] , 
        \sr_new[5] , \sr_new[4] , \sr_new[3] , \sr_new[2] , 
        \sr_new[1] , \sr_new[0] }), .sr_new_0_0(\sr_new_0[12] ), 
        .integral_0_0(\integral_0[25] ), .integral_1_0(
        \integral_1[25] ), .sum_39(\sum[39] ), .sum_14(\sum[14] ), 
        .sum_20(\sum[20] ), .sum_19(\sum[19] ), .sum_22(\sum[22] ), 
        .sum_13(\sum[13] ), .sum_17(\sum[17] ), .sum_18(\sum[18] ), 
        .sum_23(\sum[23] ), .sum_21(\sum[21] ), .sum_16(\sum[16] ), 
        .sum_15(\sum[15] ), .sum_12(\sum[12] ), .sum_11(\sum[11] ), 
        .sum_6(\sum[6] ), .sum_9(\sum[9] ), .sum_10(\sum[10] ), .sum_5(
        \sum[5] ), .sum_8(\sum[8] ), .sum_7(\sum[7] ), .sum_4(\sum[4] )
        , .sum_2_d0(\sum[2] ), .sum_1_d0(\sum[1] ), .sum_0_d0(\sum[0] )
        , .sum_3(\sum[3] ), .sum_0_0(\sum_0[39] ), .sum_1_0(
        \sum_1[39] ), .sum_2_0(\sum_2[39] ), .sum_enable(sum_enable), 
        .sum_rdy(sum_rdy), .n_rst_c(n_rst_c), .clk_c(clk_c));
    sig_gen_7 VD_SIG (.vd_done(vd_done), .n_rst_c(n_rst_c), .clk_c(
        clk_c), .sig_old_i_0(sig_old_i_0_0), .sig_prev(sig_prev_0));
    spi_rx_12s_3_1 SPI (.cur_vd({\cur_vd[11] , \cur_vd[10] , 
        \cur_vd[9] , \cur_vd[8] , \cur_vd[7] , \cur_vd[6] , 
        \cur_vd[5] , \cur_vd[4] , \cur_vd[3] , \cur_vd[2] , 
        \cur_vd[1] , \cur_vd[0] }), .vd_done(vd_done), .cs_i_1_i(
        cs_i_1_i), .sck_5_c(sck_5_c), .n_rst_c(n_rst_c), .din_15_c(
        din_15_c));
    integral_calc_13s_0_4_3 INTCALC (.sr_new({\sr_new[12] , 
        \sr_new[11] , \sr_new[10] , \sr_new[9] , \sr_new[8] , 
        \sr_new[7] , \sr_new[6] , \sr_new[5] , \sr_new[4] , 
        \sr_new[3] , \sr_new[2] , \sr_new[1] , \sr_new[0] }), .sr_old({
        \sr_old[12] , \sr_old[11] , \sr_old[10] , \sr_old[9] , 
        \sr_old[8] , \sr_old[7] , \sr_old[6] , \sr_old[5] , 
        \sr_old[4] , \sr_old[3] , \sr_old[2] , \sr_old[1] , 
        \sr_old[0] }), .sr_new_0_0(\sr_new_0[12] ), .integral({
        \integral[25] , \integral[24] , \integral[23] , \integral[22] , 
        \integral[21] , \integral[20] , \integral[19] , \integral[18] , 
        \integral[17] , \integral[16] , \integral[15] , \integral[14] , 
        \integral[13] , \integral[12] , \integral[11] , \integral[10] , 
        \integral[9] , \integral[8] , \integral[7] , \integral[6] }), 
        .integral_i({\integral_i[25] , \integral_i[24] }), 
        .integral_0_0(\integral_0[25] ), .integral_1_0(
        \integral_1[25] ), .calc_int(calc_int), .N_46_1(N_46_1_0), 
        .n_rst_c(n_rst_c), .clk_c(clk_c));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    error_calc_13s_12s_4_3 EC (.cur_error({\cur_error[12] , 
        \cur_error[11] , \cur_error[10] , \cur_error[9] , 
        \cur_error[8] , \cur_error[7] , \cur_error[6] , \cur_error[5] , 
        \cur_error[4] , \cur_error[3] , \cur_error[2] , \cur_error[1] , 
        \cur_error[0] }), .LED_15_i_0(\LED_15_i[5] ), .LED_15({
        LED_15[7], LED_15[6], LED_15[5], LED_15[4], LED_15[3], 
        LED_15[2], LED_15[1], LED_15[0]}), .average({\average[6] , 
        \average[5] , \average[4] , \average[3] , \average[2] }), 
        .calc_error(calc_error), .n_rst_c(n_rst_c), .clk_c(clk_c));
    derivative_calc_13s_4_3 DCALC (.derivative_0(\derivative[12] ), 
        .sr_prev({\sr_prev[12] , \sr_prev[11] , \sr_prev[10] , 
        \sr_prev[9] , \sr_prev[8] , \sr_prev[7] , \sr_prev[6] , 
        \sr_prev[5] , \sr_prev[4] , \sr_prev[3] , \sr_prev[2] , 
        \sr_prev[1] , \sr_prev[0] }), .sr_new({\sr_new[12] , 
        \sr_new[11] , \sr_new[10] , \sr_new[9] , \sr_new[8] , 
        \sr_new[7] , \sr_new[6] , \sr_new[5] , \sr_new[4] , 
        \sr_new[3] , \sr_new[2] , \sr_new[1] , \sr_new[0] }), 
        .deriv_enable(deriv_enable), .n_rst_c(n_rst_c), .clk_c(clk_c));
    pwm_tx_200s_32s_13s_10_1000000s_45s PWM_TX (.off_div({
        \off_div[31] , \off_div[30] , \off_div[29] , \off_div[28] , 
        \off_div[27] , \off_div[26] , \off_div[25] , \off_div[24] , 
        \off_div[23] , \off_div[22] , \off_div[21] , \off_div[20] , 
        \off_div[19] , \off_div[18] , \off_div[17] , \off_div[16] , 
        \off_div[15] , \off_div[14] , \off_div[13] , \off_div[12] , 
        \off_div[11] , \off_div[10] , \off_div[9] , \off_div[8] , 
        \off_div[7] , \off_div[6] , \off_div[5] , \off_div[4] , 
        \off_div[3] , \off_div[2] , \off_div[1] , \off_div[0] }), 
        .act_ctl_5_0(act_ctl_5_0), .pwm_chg(pwm_chg), .pwm_chg_0(
        pwm_chg_0), .n_rst_c(n_rst_c), .clk_c(clk_c), .act_ctl_5_8(
        act_ctl_5_8), .act_ctl_5_7(act_ctl_5_7), .act_ctl_5_2(
        act_ctl_5_2), .act_ctl_5_4(act_ctl_5_4), .act_ctl_5_3(
        act_ctl_5_3), .primary_15_c(primary_15_c));
    spi_clk_11s_3_1 SPICLK (.sck_5_c(sck_5_c), .n_rst_c(n_rst_c), 
        .clk_c(clk_c));
    
endmodule


module sig_gen_10(
       dec_const_c,
       n_rst_c,
       clk_c,
       dec_constd
    );
input  dec_const_c;
input  n_rst_c;
input  clk_c;
output dec_constd;

    wire sig_prev_i, sig_prev_net_1, sig_old_i_0, GND, VCC;
    
    NOR2B sig_old_RNIOSVI (.A(sig_old_i_0), .B(sig_prev_net_1), .Y(
        dec_constd));
    VCC VCC_i (.Y(VCC));
    DFN1P0 sig_old (.D(sig_prev_i), .CLK(clk_c), .PRE(n_rst_c), .Q(
        sig_old_i_0));
    DFN1C0 sig_prev (.D(dec_const_c), .CLK(clk_c), .CLR(n_rst_c), .Q(
        sig_prev_net_1));
    INV sig_old_RNO (.A(sig_prev_net_1), .Y(sig_prev_i));
    GND GND_i (.Y(GND));
    
endmodule


module PSU_Top_Level(
       clk,
       n_rst,
       inc_const,
       dec_const,
       din_12,
       sck_12,
       cs_12,
       primary_12,
       secondary_12,
       din_33,
       sck_33,
       cs_33,
       primary_33,
       secondary_33,
       din_fb,
       sck_fb,
       cs_fb,
       primary_fb,
       secondary_fb,
       active_fb,
       din_5,
       sck_5,
       cs_5,
       primary_5,
       secondary_5,
       din_15,
       sck_15,
       cs_15,
       primary_15,
       secondary_15,
       LED
    );
input  clk;
input  n_rst;
input  inc_const;
input  dec_const;
input  din_12;
output sck_12;
output cs_12;
output primary_12;
output secondary_12;
input  din_33;
output sck_33;
output cs_33;
output primary_33;
output secondary_33;
input  din_fb;
output sck_fb;
output cs_fb;
output primary_fb;
output secondary_fb;
output active_fb;
input  din_5;
output sck_5;
output cs_5;
output primary_5;
output secondary_5;
input  din_15;
output sck_15;
output cs_15;
output primary_15;
output secondary_15;
output [7:0] LED;

    wire act_ctl_5, \LED_12[0] , \LED_12[1] , \LED_12[2] , \LED_12[3] , 
        \LED_12[4] , \LED_12[5] , \LED_33[0] , \LED_33[2] , 
        \LED_33[4] , \LED_33[5] , \LED_33[6] , \LED_33[7] , 
        \LED_FB[0] , \LED_FB[1] , \LED_FB[2] , \LED_FB[3] , 
        \LED_FB[5] , \LED_FB[6] , \LED_FB[7] , \LED_5[1] , \LED_5[4] , 
        \LED_5[6] , \LED_5[7] , \LED_15[0] , \LED_15[1] , \LED_15[2] , 
        \LED_15[3] , \LED_15[4] , \LED_15[5] , \LED_15[6] , 
        \LED_15[7] , \choose[0]_net_1 , \choose[1]_net_1 , 
        \choose[2]_net_1 , choose_n1, choose_n2, VCC, choose_n0, clk_c, 
        n_rst_c, inc_const_c, dec_const_c, din_12_c, cur_clk, 
        primary_12_c, din_33_c, sck_12_c, primary_33_c, din_fb_c, 
        sck_33_c, primary_fb_c, din_5_c, sck_fb_c, primary_5_c, 
        din_15_c, sck_5_c, primary_15_c, GND, \LED_c[0] , \LED_c[1] , 
        \LED_c[2] , \LED_c[3] , \LED_c[4] , \LED_c[5] , \LED_c[6] , 
        \LED_c[7] , inc_constd, dec_constd, N_45, 
        \PID_12.SPI.cs_i_1_i , \PID_33.SPI.cs_i_1_i , 
        \PID_FB.SPI.cs_i_1_i , \PID_5.SPI.cs_i_1_i , 
        \PID_15.SPI.cs_i_1_i , act_ctl_5_i, \choose_0[2]_net_1 , 
        act_ctl_5_0, act_ctl_5_1, act_ctl_5_2, act_ctl_5_3, 
        act_ctl_5_4, act_ctl_5_5, act_ctl_5_6, act_ctl_5_7, 
        act_ctl_5_8, act_ctl_5_9;
    
    OUTBUF sck_fb_pad (.D(sck_33_c), .PAD(sck_fb));
    DFN1C0 \choose_0[2]  (.D(choose_n2), .CLK(clk_c), .CLR(n_rst_c), 
        .Q(\choose_0[2]_net_1 ));
    INBUF din_15_pad (.PAD(din_15), .Y(din_15_c));
    OUTBUF secondary_12_pad (.D(GND), .PAD(secondary_12));
    DFN1C0 \choose[1]  (.D(choose_n1), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \choose[1]_net_1 ));
    OUTBUF secondary_5_pad (.D(GND), .PAD(secondary_5));
    OUTBUF secondary_33_pad (.D(GND), .PAD(secondary_33));
    OUTBUF primary_fb_pad (.D(primary_fb_c), .PAD(primary_fb));
    sig_gen_9 INC_SIG (.inc_const_c(inc_const_c), .n_rst_c(n_rst_c), 
        .clk_c(clk_c), .inc_constd(inc_constd));
    OUTBUF sck_15_pad (.D(sck_5_c), .PAD(sck_15));
    OUTBUF cs_12_pad (.D(\PID_12.SPI.cs_i_1_i ), .PAD(cs_12));
    OUTBUF secondary_fb_pad (.D(GND), .PAD(secondary_fb));
    VCC VCC_i (.Y(VCC));
    CLKBUF n_rst_pad (.PAD(n_rst), .Y(n_rst_c));
    INBUF inc_const_pad (.PAD(inc_const), .Y(inc_const_c));
    OUTBUF \LED_pad[3]  (.D(\LED_c[3] ), .PAD(LED[3]));
    OUTBUF sck_33_pad (.D(sck_12_c), .PAD(sck_33));
    OUTBUF cs_5_pad (.D(\PID_5.SPI.cs_i_1_i ), .PAD(cs_5));
    OUTBUF \LED_pad[6]  (.D(\LED_c[6] ), .PAD(LED[6]));
    OUTBUF cs_33_pad (.D(\PID_33.SPI.cs_i_1_i ), .PAD(cs_33));
    OUTBUF \LED_pad[5]  (.D(\LED_c[5] ), .PAD(LED[5]));
    OUTBUF sck_12_pad (.D(cur_clk), .PAD(sck_12));
    OUTBUF primary_15_pad (.D(primary_15_c), .PAD(primary_15));
    OUTBUF sck_5_pad (.D(sck_fb_c), .PAD(sck_5));
    PID_controller_Z3_0 PID_FB (.LED_12_0(\LED_12[4] ), .LED_15_0(
        \LED_15[4] ), .choose_0_0(\choose_0[2]_net_1 ), .LED_c_0(
        \LED_c[4] ), .LED_5_0(\LED_5[4] ), .choose({\choose[2]_net_1 , 
        \choose[1]_net_1 , \choose[0]_net_1 }), .LED_33_0(\LED_33[4] ), 
        .LED_FB({\LED_FB[7] , \LED_FB[6] , \LED_FB[5] , nc0, 
        \LED_FB[3] , \LED_FB[2] , \LED_FB[1] , \LED_FB[0] }), 
        .primary_fb_c(primary_fb_c), .act_ctl_5(act_ctl_5), 
        .act_ctl_5_8(act_ctl_5_8), .act_ctl_5_9(act_ctl_5_9), 
        .act_ctl_5_1(act_ctl_5_1), .act_ctl_5_2(act_ctl_5_2), 
        .act_ctl_5_0(act_ctl_5_0), .act_ctl_5_3(act_ctl_5_3), 
        .act_ctl_5_i(act_ctl_5_i), .din_fb_c(din_fb_c), .cs_i_1_i(
        \PID_FB.SPI.cs_i_1_i ), .sck_33_c(sck_33_c), .clk_c(clk_c), 
        .n_rst_c(n_rst_c));
    OUTBUF \LED_pad[4]  (.D(\LED_c[4] ), .PAD(LED[4]));
    OUTBUF primary_12_pad (.D(primary_12_c), .PAD(primary_12));
    DFN1C0 \choose[0]  (.D(choose_n0), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \choose[0]_net_1 ));
    INBUF din_33_pad (.PAD(din_33), .Y(din_33_c));
    PSU_controller PSU_CTL (.act_ctl_5(act_ctl_5), .act_ctl_5_i(
        act_ctl_5_i), .act_ctl_5_0(act_ctl_5_0), .act_ctl_5_1(
        act_ctl_5_1), .act_ctl_5_2(act_ctl_5_2), .act_ctl_5_3(
        act_ctl_5_3), .act_ctl_5_4(act_ctl_5_4), .act_ctl_5_5(
        act_ctl_5_5), .act_ctl_5_6(act_ctl_5_6), .act_ctl_5_7(
        act_ctl_5_7), .act_ctl_5_8(act_ctl_5_8), .n_rst_c(n_rst_c), 
        .clk_c(clk_c), .act_ctl_5_9(act_ctl_5_9));
    GND GND_i (.Y(GND));
    OUTBUF secondary_15_pad (.D(GND), .PAD(secondary_15));
    OUTBUF \LED_pad[1]  (.D(\LED_c[1] ), .PAD(LED[1]));
    PID_controller_Z3_1 PID_33 (.choose_0_0(\choose_0[2]_net_1 ), 
        .choose({\choose[2]_net_1 , \choose[1]_net_1 , 
        \choose[0]_net_1 }), .LED_FB_2(\LED_FB[3] ), .LED_FB_0(
        \LED_FB[1] ), .LED_5_0(\LED_5[1] ), .LED_c_2(\LED_c[3] ), 
        .LED_c_0(\LED_c[1] ), .LED_12_0(\LED_12[1] ), .LED_15_0(
        \LED_15[1] ), .LED_33_0(\LED_33[0] ), .LED_33_2(\LED_33[2] ), 
        .LED_33_4(\LED_33[4] ), .LED_33_5(\LED_33[5] ), .LED_33_6(
        \LED_33[6] ), .LED_33_7(\LED_33[7] ), .primary_33_c(
        primary_33_c), .act_ctl_5(act_ctl_5), .act_ctl_5_4(act_ctl_5_4)
        , .act_ctl_5_5(act_ctl_5_5), .act_ctl_5_6(act_ctl_5_6), 
        .act_ctl_5_0(act_ctl_5_0), .act_ctl_5_3(act_ctl_5_3), 
        .act_ctl_5_1(act_ctl_5_1), .act_ctl_5_i(act_ctl_5_i), 
        .din_33_c(din_33_c), .cs_i_1_i(\PID_33.SPI.cs_i_1_i ), 
        .sck_12_c(sck_12_c), .choose_n2(choose_n2), .inc_constd(
        inc_constd), .choose_n1(choose_n1), .N_45(N_45), .dec_constd(
        dec_constd), .choose_n0(choose_n0), .clk_c(clk_c), .n_rst_c(
        n_rst_c));
    INBUF din_12_pad (.PAD(din_12), .Y(din_12_c));
    OUTBUF \LED_pad[0]  (.D(\LED_c[0] ), .PAD(LED[0]));
    INBUF dec_const_pad (.PAD(dec_const), .Y(dec_const_c));
    PID_controller_Z4 PID_5 (.choose_0_0(\choose_0[2]_net_1 ), 
        .LED_12_0(\LED_12[0] ), .LED_12_2(\LED_12[2] ), .LED_12_3(
        \LED_12[3] ), .LED_12_5(\LED_12[5] ), .LED_15_0(\LED_15[0] ), 
        .LED_15_2(\LED_15[2] ), .LED_15_3(\LED_15[3] ), .LED_15_5(
        \LED_15[5] ), .LED_c_0(\LED_c[0] ), .LED_c_2(\LED_c[2] ), 
        .LED_c_5(\LED_c[5] ), .choose({\choose[2]_net_1 , 
        \choose[1]_net_1 , \choose[0]_net_1 }), .LED_FB_0(\LED_FB[0] ), 
        .LED_FB_2(\LED_FB[2] ), .LED_FB_5(\LED_FB[5] ), .LED_33_0(
        \LED_33[0] ), .LED_33_2(\LED_33[2] ), .LED_33_5(\LED_33[5] ), 
        .LED_5_0(\LED_5[1] ), .LED_5_3(\LED_5[4] ), .LED_5_5(
        \LED_5[6] ), .LED_5_6(\LED_5[7] ), .primary_5_c(primary_5_c), 
        .act_ctl_5_4(act_ctl_5_4), .act_ctl_5_8(act_ctl_5_8), 
        .act_ctl_5_6(act_ctl_5_6), .act_ctl_5_7(act_ctl_5_7), 
        .act_ctl_5_0(act_ctl_5_0), .act_ctl_5_1(act_ctl_5_1), 
        .act_ctl_5_i(act_ctl_5_i), .N_45(N_45), .din_5_c(din_5_c), 
        .cs_i_1_i(\PID_5.SPI.cs_i_1_i ), .sck_fb_c(sck_fb_c), .clk_c(
        clk_c), .n_rst_c(n_rst_c));
    PID_controller_Z2 PID_12 (.choose_0_0(\choose_0[2]_net_1 ), 
        .choose({\choose[2]_net_1 , \choose[1]_net_1 , 
        \choose[0]_net_1 }), .LED_15({\LED_15[7] , \LED_15[6] }), 
        .LED_c({\LED_c[7] , \LED_c[6] }), .LED_5({\LED_5[7] , 
        \LED_5[6] }), .LED_FB({\LED_FB[7] , \LED_FB[6] }), .LED_33({
        \LED_33[7] , \LED_33[6] }), .LED_12({\LED_12[5] , \LED_12[4] , 
        \LED_12[3] , \LED_12[2] , \LED_12[1] , \LED_12[0] }), 
        .primary_12_c(primary_12_c), .act_ctl_5_7(act_ctl_5_7), 
        .act_ctl_5_3(act_ctl_5_3), .act_ctl_5_4(act_ctl_5_4), 
        .act_ctl_5_9(act_ctl_5_9), .act_ctl_5(act_ctl_5), .act_ctl_5_8(
        act_ctl_5_8), .act_ctl_5_0(act_ctl_5_0), .act_ctl_5_i(
        act_ctl_5_i), .din_12_c(din_12_c), .cs_i_1_i(
        \PID_12.SPI.cs_i_1_i ), .cur_clk(cur_clk), .clk_c(clk_c), 
        .n_rst_c(n_rst_c));
    PID_controller_Z5 PID_15 (.LED_15({\LED_15[7] , \LED_15[6] , 
        \LED_15[5] , \LED_15[4] , \LED_15[3] , \LED_15[2] , 
        \LED_15[1] , \LED_15[0] }), .primary_15_c(primary_15_c), 
        .act_ctl_5_3(act_ctl_5_3), .act_ctl_5_4(act_ctl_5_4), 
        .act_ctl_5_2(act_ctl_5_2), .act_ctl_5_7(act_ctl_5_7), 
        .act_ctl_5_8(act_ctl_5_8), .act_ctl_5_0(act_ctl_5_0), 
        .din_15_c(din_15_c), .cs_i_1_i(\PID_15.SPI.cs_i_1_i ), 
        .sck_5_c(sck_5_c), .clk_c(clk_c), .n_rst_c(n_rst_c));
    OUTBUF primary_33_pad (.D(primary_33_c), .PAD(primary_33));
    OUTBUF \LED_pad[7]  (.D(\LED_c[7] ), .PAD(LED[7]));
    OUTBUF primary_5_pad (.D(primary_5_c), .PAD(primary_5));
    DFN1C0 \choose[2]  (.D(choose_n2), .CLK(clk_c), .CLR(n_rst_c), .Q(
        \choose[2]_net_1 ));
    OUTBUF active_fb_pad (.D(GND), .PAD(active_fb));
    OUTBUF cs_fb_pad (.D(\PID_FB.SPI.cs_i_1_i ), .PAD(cs_fb));
    OUTBUF cs_15_pad (.D(\PID_15.SPI.cs_i_1_i ), .PAD(cs_15));
    OUTBUF \LED_pad[2]  (.D(\LED_c[2] ), .PAD(LED[2]));
    sig_gen_10 DEC_SIG (.dec_const_c(dec_const_c), .n_rst_c(n_rst_c), 
        .clk_c(clk_c), .dec_constd(dec_constd));
    INBUF din_5_pad (.PAD(din_5), .Y(din_5_c));
    INBUF din_fb_pad (.PAD(din_fb), .Y(din_fb_c));
    CLKBUF clk_pad (.PAD(clk), .Y(clk_c));
    
endmodule
