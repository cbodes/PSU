///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: error_calc.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::ProASIC3E> <Die::A3PE1500> <Package::208 PQFP>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

//`timescale <time_units> / <precision>

module error_calc #(
    parameter ADC_WIDTH = 8,
    parameter SPI_WIDTH = 13
) (   
    input clk, n_rst, calc_error,
    input [ADC_WIDTH-1:0] target_v,
    input [ADC_WIDTH-1:0] cur_vd,
    output reg [ADC_WIDTH-1:0] diff
);
    
reg [ADC_WIDTH-1:0] diffreg;

//assign diff = {diffreg[ADC_WIDTH-1], 2'b00, diffreg[ADC_WIDTH-2:2]};
assign diff = diffreg;

always @(posedge clk, negedge n_rst) begin
    if (n_rst == 0) begin
        diffreg <= '0;
    end else if (calc_error == 1) begin
        diffreg <= cur_vd - target_v;
    end
end

endmodule

